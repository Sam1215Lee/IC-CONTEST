
module lcd_ctrl ( clk, reset, datain, cmd, cmd_valid, dataout, output_valid, 
        busy );
  input [7:0] datain;
  input [2:0] cmd;
  output [7:0] dataout;
  input clk, reset, cmd_valid;
  output output_valid, busy;
  wire   next, N198, N199, N200, N201, \col_t[2] , N449, N450, N451, N452, n78,
         n84, n85, n86, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, \add_0_root_add_171_2/carry[5] ,
         \add_0_root_add_171_2/carry[3] , \add_0_root_add_171_2/carry[2] ,
         \add_1_root_add_171_2/carry[4] , \add_1_root_add_171_2/carry[3] ,
         \r407/carry[5] , \r407/carry[4] , \r407/carry[3] , \r407/carry[2] ,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090;
  wire   [5:0] cnt;
  wire   [2:0] row;
  wire   [5:0] outpos;
  wire   [2:0] row_t;

  DFFRXL \cnt_reg[5]  ( .D(n740), .CK(clk), .RN(n1054), .Q(n745), .QN(n91) );
  DFFRXL cur_reg ( .D(next), .CK(clk), .RN(n1054), .Q(n744), .QN(n78) );
  DFFRXL \cmdreg_reg[1]  ( .D(n737), .CK(clk), .RN(n1054), .Q(n747), .QN(n85)
         );
  DFFRXL \cmdreg_reg[0]  ( .D(n738), .CK(clk), .RN(n1054), .Q(n743), .QN(n86)
         );
  DFFRXL \cmdreg_reg[2]  ( .D(n739), .CK(clk), .RN(n1054), .Q(n742), .QN(n84)
         );
  EDFFX1 \data_reg[0][7]  ( .D(datain[7]), .E(n1055), .CK(clk), .QN(n97) );
  EDFFX1 \data_reg[0][6]  ( .D(datain[6]), .E(n1055), .CK(clk), .QN(n98) );
  EDFFX1 \data_reg[0][5]  ( .D(datain[5]), .E(n1055), .CK(clk), .QN(n99) );
  EDFFX1 \data_reg[0][4]  ( .D(datain[4]), .E(n1055), .CK(clk), .QN(n100) );
  EDFFX1 \data_reg[0][3]  ( .D(datain[3]), .E(n1055), .CK(clk), .QN(n101) );
  EDFFX1 \data_reg[0][2]  ( .D(datain[2]), .E(n1055), .CK(clk), .QN(n102) );
  EDFFX1 \data_reg[0][1]  ( .D(datain[1]), .E(n1055), .CK(clk), .QN(n103) );
  EDFFX1 \data_reg[0][0]  ( .D(datain[0]), .E(n1055), .CK(clk), .QN(n104) );
  EDFFX1 \data_reg[1][7]  ( .D(datain[7]), .E(n1056), .CK(clk), .QN(n105) );
  EDFFX1 \data_reg[1][6]  ( .D(datain[6]), .E(n1056), .CK(clk), .QN(n106) );
  EDFFX1 \data_reg[1][5]  ( .D(datain[5]), .E(n1056), .CK(clk), .QN(n107) );
  EDFFX1 \data_reg[1][4]  ( .D(datain[4]), .E(n1056), .CK(clk), .QN(n108) );
  EDFFX1 \data_reg[1][3]  ( .D(datain[3]), .E(n1056), .CK(clk), .QN(n109) );
  EDFFX1 \data_reg[1][2]  ( .D(datain[2]), .E(n1056), .CK(clk), .QN(n110) );
  EDFFX1 \data_reg[1][1]  ( .D(datain[1]), .E(n1056), .CK(clk), .QN(n111) );
  EDFFX1 \data_reg[1][0]  ( .D(datain[0]), .E(n1056), .CK(clk), .QN(n112) );
  EDFFX1 \data_reg[2][7]  ( .D(datain[7]), .E(n1057), .CK(clk), .QN(n113) );
  EDFFX1 \data_reg[2][6]  ( .D(datain[6]), .E(n1057), .CK(clk), .QN(n114) );
  EDFFX1 \data_reg[2][5]  ( .D(datain[5]), .E(n1057), .CK(clk), .QN(n115) );
  EDFFX1 \data_reg[2][4]  ( .D(datain[4]), .E(n1057), .CK(clk), .QN(n116) );
  EDFFX1 \data_reg[2][3]  ( .D(datain[3]), .E(n1057), .CK(clk), .QN(n117) );
  EDFFX1 \data_reg[2][2]  ( .D(datain[2]), .E(n1057), .CK(clk), .QN(n118) );
  EDFFX1 \data_reg[2][1]  ( .D(datain[1]), .E(n1057), .CK(clk), .QN(n119) );
  EDFFX1 \data_reg[2][0]  ( .D(datain[0]), .E(n1057), .CK(clk), .QN(n120) );
  EDFFX1 \data_reg[3][7]  ( .D(datain[7]), .E(n1058), .CK(clk), .QN(n121) );
  EDFFX1 \data_reg[3][6]  ( .D(datain[6]), .E(n1058), .CK(clk), .QN(n122) );
  EDFFX1 \data_reg[3][5]  ( .D(datain[5]), .E(n1058), .CK(clk), .QN(n123) );
  EDFFX1 \data_reg[3][4]  ( .D(datain[4]), .E(n1058), .CK(clk), .QN(n124) );
  EDFFX1 \data_reg[3][3]  ( .D(datain[3]), .E(n1058), .CK(clk), .QN(n125) );
  EDFFX1 \data_reg[3][2]  ( .D(datain[2]), .E(n1058), .CK(clk), .QN(n126) );
  EDFFX1 \data_reg[3][1]  ( .D(datain[1]), .E(n1058), .CK(clk), .QN(n127) );
  EDFFX1 \data_reg[3][0]  ( .D(datain[0]), .E(n1058), .CK(clk), .QN(n128) );
  EDFFX1 \data_reg[4][7]  ( .D(datain[7]), .E(n1059), .CK(clk), .QN(n129) );
  EDFFX1 \data_reg[4][6]  ( .D(datain[6]), .E(n1059), .CK(clk), .QN(n130) );
  EDFFX1 \data_reg[4][5]  ( .D(datain[5]), .E(n1059), .CK(clk), .QN(n131) );
  EDFFX1 \data_reg[4][4]  ( .D(datain[4]), .E(n1059), .CK(clk), .QN(n132) );
  EDFFX1 \data_reg[4][3]  ( .D(datain[3]), .E(n1059), .CK(clk), .QN(n133) );
  EDFFX1 \data_reg[4][2]  ( .D(datain[2]), .E(n1059), .CK(clk), .QN(n134) );
  EDFFX1 \data_reg[4][1]  ( .D(datain[1]), .E(n1059), .CK(clk), .QN(n135) );
  EDFFX1 \data_reg[4][0]  ( .D(datain[0]), .E(n1059), .CK(clk), .QN(n136) );
  EDFFX1 \data_reg[5][7]  ( .D(datain[7]), .E(n1060), .CK(clk), .QN(n137) );
  EDFFX1 \data_reg[5][6]  ( .D(datain[6]), .E(n1060), .CK(clk), .QN(n138) );
  EDFFX1 \data_reg[5][5]  ( .D(datain[5]), .E(n1060), .CK(clk), .QN(n139) );
  EDFFX1 \data_reg[5][4]  ( .D(datain[4]), .E(n1060), .CK(clk), .QN(n140) );
  EDFFX1 \data_reg[5][3]  ( .D(datain[3]), .E(n1060), .CK(clk), .QN(n141) );
  EDFFX1 \data_reg[5][2]  ( .D(datain[2]), .E(n1060), .CK(clk), .QN(n142) );
  EDFFX1 \data_reg[5][1]  ( .D(datain[1]), .E(n1060), .CK(clk), .QN(n143) );
  EDFFX1 \data_reg[5][0]  ( .D(datain[0]), .E(n1060), .CK(clk), .QN(n144) );
  EDFFX1 \data_reg[6][7]  ( .D(datain[7]), .E(n1061), .CK(clk), .QN(n145) );
  EDFFX1 \data_reg[6][6]  ( .D(datain[6]), .E(n1061), .CK(clk), .QN(n146) );
  EDFFX1 \data_reg[6][5]  ( .D(datain[5]), .E(n1061), .CK(clk), .QN(n147) );
  EDFFX1 \data_reg[6][4]  ( .D(datain[4]), .E(n1061), .CK(clk), .QN(n148) );
  EDFFX1 \data_reg[6][3]  ( .D(datain[3]), .E(n1061), .CK(clk), .QN(n149) );
  EDFFX1 \data_reg[6][2]  ( .D(datain[2]), .E(n1061), .CK(clk), .QN(n150) );
  EDFFX1 \data_reg[6][1]  ( .D(datain[1]), .E(n1061), .CK(clk), .QN(n151) );
  EDFFX1 \data_reg[6][0]  ( .D(datain[0]), .E(n1061), .CK(clk), .QN(n152) );
  EDFFX1 \data_reg[7][7]  ( .D(datain[7]), .E(n1062), .CK(clk), .QN(n153) );
  EDFFX1 \data_reg[7][6]  ( .D(datain[6]), .E(n1062), .CK(clk), .QN(n154) );
  EDFFX1 \data_reg[7][5]  ( .D(datain[5]), .E(n1062), .CK(clk), .QN(n155) );
  EDFFX1 \data_reg[7][4]  ( .D(datain[4]), .E(n1062), .CK(clk), .QN(n156) );
  EDFFX1 \data_reg[7][3]  ( .D(datain[3]), .E(n1062), .CK(clk), .QN(n157) );
  EDFFX1 \data_reg[7][2]  ( .D(datain[2]), .E(n1062), .CK(clk), .QN(n158) );
  EDFFX1 \data_reg[7][1]  ( .D(datain[1]), .E(n1062), .CK(clk), .QN(n159) );
  EDFFX1 \data_reg[7][0]  ( .D(datain[0]), .E(n1062), .CK(clk), .QN(n160) );
  EDFFX1 \data_reg[8][7]  ( .D(datain[7]), .E(n1063), .CK(clk), .QN(n161) );
  EDFFX1 \data_reg[8][6]  ( .D(datain[6]), .E(n1063), .CK(clk), .QN(n162) );
  EDFFX1 \data_reg[8][5]  ( .D(datain[5]), .E(n1063), .CK(clk), .QN(n163) );
  EDFFX1 \data_reg[8][4]  ( .D(datain[4]), .E(n1063), .CK(clk), .QN(n164) );
  EDFFX1 \data_reg[8][3]  ( .D(datain[3]), .E(n1063), .CK(clk), .QN(n165) );
  EDFFX1 \data_reg[8][2]  ( .D(datain[2]), .E(n1063), .CK(clk), .QN(n166) );
  EDFFX1 \data_reg[8][1]  ( .D(datain[1]), .E(n1063), .CK(clk), .QN(n167) );
  EDFFX1 \data_reg[8][0]  ( .D(datain[0]), .E(n1063), .CK(clk), .QN(n168) );
  EDFFX1 \data_reg[9][7]  ( .D(datain[7]), .E(n1064), .CK(clk), .QN(n169) );
  EDFFX1 \data_reg[9][6]  ( .D(datain[6]), .E(n1064), .CK(clk), .QN(n170) );
  EDFFX1 \data_reg[9][5]  ( .D(datain[5]), .E(n1064), .CK(clk), .QN(n171) );
  EDFFX1 \data_reg[9][4]  ( .D(datain[4]), .E(n1064), .CK(clk), .QN(n172) );
  EDFFX1 \data_reg[9][3]  ( .D(datain[3]), .E(n1064), .CK(clk), .QN(n173) );
  EDFFX1 \data_reg[9][2]  ( .D(datain[2]), .E(n1064), .CK(clk), .QN(n174) );
  EDFFX1 \data_reg[9][1]  ( .D(datain[1]), .E(n1064), .CK(clk), .QN(n175) );
  EDFFX1 \data_reg[9][0]  ( .D(datain[0]), .E(n1064), .CK(clk), .QN(n176) );
  EDFFX1 \data_reg[10][7]  ( .D(datain[7]), .E(n1065), .CK(clk), .QN(n177) );
  EDFFX1 \data_reg[10][6]  ( .D(datain[6]), .E(n1065), .CK(clk), .QN(n178) );
  EDFFX1 \data_reg[10][5]  ( .D(datain[5]), .E(n1065), .CK(clk), .QN(n179) );
  EDFFX1 \data_reg[10][4]  ( .D(datain[4]), .E(n1065), .CK(clk), .QN(n180) );
  EDFFX1 \data_reg[10][3]  ( .D(datain[3]), .E(n1065), .CK(clk), .QN(n181) );
  EDFFX1 \data_reg[10][2]  ( .D(datain[2]), .E(n1065), .CK(clk), .QN(n182) );
  EDFFX1 \data_reg[10][1]  ( .D(datain[1]), .E(n1065), .CK(clk), .QN(n183) );
  EDFFX1 \data_reg[10][0]  ( .D(datain[0]), .E(n1065), .CK(clk), .QN(n184) );
  EDFFX1 \data_reg[11][7]  ( .D(datain[7]), .E(n1066), .CK(clk), .QN(n185) );
  EDFFX1 \data_reg[11][6]  ( .D(datain[6]), .E(n1066), .CK(clk), .QN(n186) );
  EDFFX1 \data_reg[11][5]  ( .D(datain[5]), .E(n1066), .CK(clk), .QN(n187) );
  EDFFX1 \data_reg[11][4]  ( .D(datain[4]), .E(n1066), .CK(clk), .QN(n188) );
  EDFFX1 \data_reg[11][3]  ( .D(datain[3]), .E(n1066), .CK(clk), .QN(n189) );
  EDFFX1 \data_reg[11][2]  ( .D(datain[2]), .E(n1066), .CK(clk), .QN(n190) );
  EDFFX1 \data_reg[11][1]  ( .D(datain[1]), .E(n1066), .CK(clk), .QN(n191) );
  EDFFX1 \data_reg[11][0]  ( .D(datain[0]), .E(n1066), .CK(clk), .QN(n192) );
  EDFFX1 \data_reg[12][7]  ( .D(datain[7]), .E(n1067), .CK(clk), .QN(n193) );
  EDFFX1 \data_reg[12][6]  ( .D(datain[6]), .E(n1067), .CK(clk), .QN(n194) );
  EDFFX1 \data_reg[12][5]  ( .D(datain[5]), .E(n1067), .CK(clk), .QN(n195) );
  EDFFX1 \data_reg[12][4]  ( .D(datain[4]), .E(n1067), .CK(clk), .QN(n196) );
  EDFFX1 \data_reg[12][3]  ( .D(datain[3]), .E(n1067), .CK(clk), .QN(n197) );
  EDFFX1 \data_reg[12][2]  ( .D(datain[2]), .E(n1067), .CK(clk), .QN(n198) );
  EDFFX1 \data_reg[12][1]  ( .D(datain[1]), .E(n1067), .CK(clk), .QN(n199) );
  EDFFX1 \data_reg[12][0]  ( .D(datain[0]), .E(n1067), .CK(clk), .QN(n200) );
  EDFFX1 \data_reg[13][7]  ( .D(datain[7]), .E(n1068), .CK(clk), .QN(n201) );
  EDFFX1 \data_reg[13][6]  ( .D(datain[6]), .E(n1068), .CK(clk), .QN(n202) );
  EDFFX1 \data_reg[13][5]  ( .D(datain[5]), .E(n1068), .CK(clk), .QN(n203) );
  EDFFX1 \data_reg[13][4]  ( .D(datain[4]), .E(n1068), .CK(clk), .QN(n204) );
  EDFFX1 \data_reg[13][3]  ( .D(datain[3]), .E(n1068), .CK(clk), .QN(n205) );
  EDFFX1 \data_reg[13][2]  ( .D(datain[2]), .E(n1068), .CK(clk), .QN(n206) );
  EDFFX1 \data_reg[13][1]  ( .D(datain[1]), .E(n1068), .CK(clk), .QN(n207) );
  EDFFX1 \data_reg[13][0]  ( .D(datain[0]), .E(n1068), .CK(clk), .QN(n208) );
  EDFFX1 \data_reg[14][7]  ( .D(datain[7]), .E(n1069), .CK(clk), .QN(n209) );
  EDFFX1 \data_reg[14][6]  ( .D(datain[6]), .E(n1069), .CK(clk), .QN(n210) );
  EDFFX1 \data_reg[14][5]  ( .D(datain[5]), .E(n1069), .CK(clk), .QN(n211) );
  EDFFX1 \data_reg[14][4]  ( .D(datain[4]), .E(n1069), .CK(clk), .QN(n212) );
  EDFFX1 \data_reg[14][3]  ( .D(datain[3]), .E(n1069), .CK(clk), .QN(n213) );
  EDFFX1 \data_reg[14][2]  ( .D(datain[2]), .E(n1069), .CK(clk), .QN(n214) );
  EDFFX1 \data_reg[14][1]  ( .D(datain[1]), .E(n1069), .CK(clk), .QN(n215) );
  EDFFX1 \data_reg[14][0]  ( .D(datain[0]), .E(n1069), .CK(clk), .QN(n216) );
  EDFFX1 \data_reg[15][7]  ( .D(datain[7]), .E(n1070), .CK(clk), .QN(n217) );
  EDFFX1 \data_reg[15][6]  ( .D(datain[6]), .E(n1070), .CK(clk), .QN(n218) );
  EDFFX1 \data_reg[15][5]  ( .D(datain[5]), .E(n1070), .CK(clk), .QN(n219) );
  EDFFX1 \data_reg[15][4]  ( .D(datain[4]), .E(n1070), .CK(clk), .QN(n220) );
  EDFFX1 \data_reg[15][3]  ( .D(datain[3]), .E(n1070), .CK(clk), .QN(n221) );
  EDFFX1 \data_reg[15][2]  ( .D(datain[2]), .E(n1070), .CK(clk), .QN(n222) );
  EDFFX1 \data_reg[15][1]  ( .D(datain[1]), .E(n1070), .CK(clk), .QN(n223) );
  EDFFX1 \data_reg[15][0]  ( .D(datain[0]), .E(n1070), .CK(clk), .QN(n224) );
  EDFFX1 \data_reg[16][7]  ( .D(datain[7]), .E(n1071), .CK(clk), .QN(n225) );
  EDFFX1 \data_reg[16][6]  ( .D(datain[6]), .E(n1071), .CK(clk), .QN(n226) );
  EDFFX1 \data_reg[16][5]  ( .D(datain[5]), .E(n1071), .CK(clk), .QN(n227) );
  EDFFX1 \data_reg[16][4]  ( .D(datain[4]), .E(n1071), .CK(clk), .QN(n228) );
  EDFFX1 \data_reg[16][3]  ( .D(datain[3]), .E(n1071), .CK(clk), .QN(n229) );
  EDFFX1 \data_reg[16][2]  ( .D(datain[2]), .E(n1071), .CK(clk), .QN(n230) );
  EDFFX1 \data_reg[16][1]  ( .D(datain[1]), .E(n1071), .CK(clk), .QN(n231) );
  EDFFX1 \data_reg[16][0]  ( .D(datain[0]), .E(n1071), .CK(clk), .QN(n232) );
  EDFFX1 \data_reg[17][7]  ( .D(datain[7]), .E(n1072), .CK(clk), .QN(n233) );
  EDFFX1 \data_reg[17][6]  ( .D(datain[6]), .E(n1072), .CK(clk), .QN(n234) );
  EDFFX1 \data_reg[17][5]  ( .D(datain[5]), .E(n1072), .CK(clk), .QN(n235) );
  EDFFX1 \data_reg[17][4]  ( .D(datain[4]), .E(n1072), .CK(clk), .QN(n236) );
  EDFFX1 \data_reg[17][3]  ( .D(datain[3]), .E(n1072), .CK(clk), .QN(n237) );
  EDFFX1 \data_reg[17][2]  ( .D(datain[2]), .E(n1072), .CK(clk), .QN(n238) );
  EDFFX1 \data_reg[17][1]  ( .D(datain[1]), .E(n1072), .CK(clk), .QN(n239) );
  EDFFX1 \data_reg[17][0]  ( .D(datain[0]), .E(n1072), .CK(clk), .QN(n240) );
  EDFFX1 \data_reg[18][7]  ( .D(datain[7]), .E(n1073), .CK(clk), .QN(n241) );
  EDFFX1 \data_reg[18][6]  ( .D(datain[6]), .E(n1073), .CK(clk), .QN(n242) );
  EDFFX1 \data_reg[18][5]  ( .D(datain[5]), .E(n1073), .CK(clk), .QN(n243) );
  EDFFX1 \data_reg[18][4]  ( .D(datain[4]), .E(n1073), .CK(clk), .QN(n244) );
  EDFFX1 \data_reg[18][3]  ( .D(datain[3]), .E(n1073), .CK(clk), .QN(n245) );
  EDFFX1 \data_reg[18][2]  ( .D(datain[2]), .E(n1073), .CK(clk), .QN(n246) );
  EDFFX1 \data_reg[18][1]  ( .D(datain[1]), .E(n1073), .CK(clk), .QN(n247) );
  EDFFX1 \data_reg[18][0]  ( .D(datain[0]), .E(n1073), .CK(clk), .QN(n248) );
  EDFFX1 \data_reg[19][7]  ( .D(datain[7]), .E(n1074), .CK(clk), .QN(n249) );
  EDFFX1 \data_reg[19][6]  ( .D(datain[6]), .E(n1074), .CK(clk), .QN(n250) );
  EDFFX1 \data_reg[19][5]  ( .D(datain[5]), .E(n1074), .CK(clk), .QN(n251) );
  EDFFX1 \data_reg[19][4]  ( .D(datain[4]), .E(n1074), .CK(clk), .QN(n252) );
  EDFFX1 \data_reg[19][3]  ( .D(datain[3]), .E(n1074), .CK(clk), .QN(n253) );
  EDFFX1 \data_reg[19][2]  ( .D(datain[2]), .E(n1074), .CK(clk), .QN(n254) );
  EDFFX1 \data_reg[19][1]  ( .D(datain[1]), .E(n1074), .CK(clk), .QN(n255) );
  EDFFX1 \data_reg[19][0]  ( .D(datain[0]), .E(n1074), .CK(clk), .QN(n256) );
  EDFFX1 \data_reg[20][7]  ( .D(datain[7]), .E(n1075), .CK(clk), .QN(n257) );
  EDFFX1 \data_reg[20][6]  ( .D(datain[6]), .E(n1075), .CK(clk), .QN(n258) );
  EDFFX1 \data_reg[20][5]  ( .D(datain[5]), .E(n1075), .CK(clk), .QN(n259) );
  EDFFX1 \data_reg[20][4]  ( .D(datain[4]), .E(n1075), .CK(clk), .QN(n260) );
  EDFFX1 \data_reg[20][3]  ( .D(datain[3]), .E(n1075), .CK(clk), .QN(n261) );
  EDFFX1 \data_reg[20][2]  ( .D(datain[2]), .E(n1075), .CK(clk), .QN(n262) );
  EDFFX1 \data_reg[20][1]  ( .D(datain[1]), .E(n1075), .CK(clk), .QN(n263) );
  EDFFX1 \data_reg[20][0]  ( .D(datain[0]), .E(n1075), .CK(clk), .QN(n264) );
  EDFFX1 \data_reg[21][7]  ( .D(datain[7]), .E(n1076), .CK(clk), .QN(n265) );
  EDFFX1 \data_reg[21][6]  ( .D(datain[6]), .E(n1076), .CK(clk), .QN(n266) );
  EDFFX1 \data_reg[21][5]  ( .D(datain[5]), .E(n1076), .CK(clk), .QN(n267) );
  EDFFX1 \data_reg[21][4]  ( .D(datain[4]), .E(n1076), .CK(clk), .QN(n268) );
  EDFFX1 \data_reg[21][3]  ( .D(datain[3]), .E(n1076), .CK(clk), .QN(n269) );
  EDFFX1 \data_reg[21][2]  ( .D(datain[2]), .E(n1076), .CK(clk), .QN(n270) );
  EDFFX1 \data_reg[21][1]  ( .D(datain[1]), .E(n1076), .CK(clk), .QN(n271) );
  EDFFX1 \data_reg[21][0]  ( .D(datain[0]), .E(n1076), .CK(clk), .QN(n272) );
  EDFFX1 \data_reg[22][7]  ( .D(datain[7]), .E(n1077), .CK(clk), .QN(n273) );
  EDFFX1 \data_reg[22][6]  ( .D(datain[6]), .E(n1077), .CK(clk), .QN(n274) );
  EDFFX1 \data_reg[22][5]  ( .D(datain[5]), .E(n1077), .CK(clk), .QN(n275) );
  EDFFX1 \data_reg[22][4]  ( .D(datain[4]), .E(n1077), .CK(clk), .QN(n276) );
  EDFFX1 \data_reg[22][3]  ( .D(datain[3]), .E(n1077), .CK(clk), .QN(n277) );
  EDFFX1 \data_reg[22][2]  ( .D(datain[2]), .E(n1077), .CK(clk), .QN(n278) );
  EDFFX1 \data_reg[22][1]  ( .D(datain[1]), .E(n1077), .CK(clk), .QN(n279) );
  EDFFX1 \data_reg[22][0]  ( .D(datain[0]), .E(n1077), .CK(clk), .QN(n280) );
  EDFFX1 \data_reg[23][7]  ( .D(datain[7]), .E(n1078), .CK(clk), .QN(n281) );
  EDFFX1 \data_reg[23][6]  ( .D(datain[6]), .E(n1078), .CK(clk), .QN(n282) );
  EDFFX1 \data_reg[23][5]  ( .D(datain[5]), .E(n1078), .CK(clk), .QN(n283) );
  EDFFX1 \data_reg[23][4]  ( .D(datain[4]), .E(n1078), .CK(clk), .QN(n284) );
  EDFFX1 \data_reg[23][3]  ( .D(datain[3]), .E(n1078), .CK(clk), .QN(n285) );
  EDFFX1 \data_reg[23][2]  ( .D(datain[2]), .E(n1078), .CK(clk), .QN(n286) );
  EDFFX1 \data_reg[23][1]  ( .D(datain[1]), .E(n1078), .CK(clk), .QN(n287) );
  EDFFX1 \data_reg[23][0]  ( .D(datain[0]), .E(n1078), .CK(clk), .QN(n288) );
  EDFFX1 \data_reg[24][7]  ( .D(datain[7]), .E(n1079), .CK(clk), .QN(n289) );
  EDFFX1 \data_reg[24][6]  ( .D(datain[6]), .E(n1079), .CK(clk), .QN(n290) );
  EDFFX1 \data_reg[24][5]  ( .D(datain[5]), .E(n1079), .CK(clk), .QN(n291) );
  EDFFX1 \data_reg[24][4]  ( .D(datain[4]), .E(n1079), .CK(clk), .QN(n292) );
  EDFFX1 \data_reg[24][3]  ( .D(datain[3]), .E(n1079), .CK(clk), .QN(n293) );
  EDFFX1 \data_reg[24][2]  ( .D(datain[2]), .E(n1079), .CK(clk), .QN(n294) );
  EDFFX1 \data_reg[24][1]  ( .D(datain[1]), .E(n1079), .CK(clk), .QN(n295) );
  EDFFX1 \data_reg[24][0]  ( .D(datain[0]), .E(n1079), .CK(clk), .QN(n296) );
  EDFFX1 \data_reg[25][7]  ( .D(datain[7]), .E(n1080), .CK(clk), .QN(n297) );
  EDFFX1 \data_reg[25][6]  ( .D(datain[6]), .E(n1080), .CK(clk), .QN(n298) );
  EDFFX1 \data_reg[25][5]  ( .D(datain[5]), .E(n1080), .CK(clk), .QN(n299) );
  EDFFX1 \data_reg[25][4]  ( .D(datain[4]), .E(n1080), .CK(clk), .QN(n300) );
  EDFFX1 \data_reg[25][3]  ( .D(datain[3]), .E(n1080), .CK(clk), .QN(n301) );
  EDFFX1 \data_reg[25][2]  ( .D(datain[2]), .E(n1080), .CK(clk), .QN(n302) );
  EDFFX1 \data_reg[25][1]  ( .D(datain[1]), .E(n1080), .CK(clk), .QN(n303) );
  EDFFX1 \data_reg[25][0]  ( .D(datain[0]), .E(n1080), .CK(clk), .QN(n304) );
  EDFFX1 \data_reg[26][7]  ( .D(datain[7]), .E(n1081), .CK(clk), .QN(n305) );
  EDFFX1 \data_reg[26][6]  ( .D(datain[6]), .E(n1081), .CK(clk), .QN(n306) );
  EDFFX1 \data_reg[26][5]  ( .D(datain[5]), .E(n1081), .CK(clk), .QN(n307) );
  EDFFX1 \data_reg[26][4]  ( .D(datain[4]), .E(n1081), .CK(clk), .QN(n308) );
  EDFFX1 \data_reg[26][3]  ( .D(datain[3]), .E(n1081), .CK(clk), .QN(n309) );
  EDFFX1 \data_reg[26][2]  ( .D(datain[2]), .E(n1081), .CK(clk), .QN(n310) );
  EDFFX1 \data_reg[26][1]  ( .D(datain[1]), .E(n1081), .CK(clk), .QN(n311) );
  EDFFX1 \data_reg[26][0]  ( .D(datain[0]), .E(n1081), .CK(clk), .QN(n312) );
  EDFFX1 \data_reg[27][7]  ( .D(datain[7]), .E(n1082), .CK(clk), .QN(n313) );
  EDFFX1 \data_reg[27][6]  ( .D(datain[6]), .E(n1082), .CK(clk), .QN(n314) );
  EDFFX1 \data_reg[27][5]  ( .D(datain[5]), .E(n1082), .CK(clk), .QN(n315) );
  EDFFX1 \data_reg[27][4]  ( .D(datain[4]), .E(n1082), .CK(clk), .QN(n316) );
  EDFFX1 \data_reg[27][3]  ( .D(datain[3]), .E(n1082), .CK(clk), .QN(n317) );
  EDFFX1 \data_reg[27][2]  ( .D(datain[2]), .E(n1082), .CK(clk), .QN(n318) );
  EDFFX1 \data_reg[27][1]  ( .D(datain[1]), .E(n1082), .CK(clk), .QN(n319) );
  EDFFX1 \data_reg[27][0]  ( .D(datain[0]), .E(n1082), .CK(clk), .QN(n320) );
  EDFFX1 \data_reg[28][7]  ( .D(datain[7]), .E(n1083), .CK(clk), .QN(n321) );
  EDFFX1 \data_reg[28][6]  ( .D(datain[6]), .E(n1083), .CK(clk), .QN(n322) );
  EDFFX1 \data_reg[28][5]  ( .D(datain[5]), .E(n1083), .CK(clk), .QN(n323) );
  EDFFX1 \data_reg[28][4]  ( .D(datain[4]), .E(n1083), .CK(clk), .QN(n324) );
  EDFFX1 \data_reg[28][3]  ( .D(datain[3]), .E(n1083), .CK(clk), .QN(n325) );
  EDFFX1 \data_reg[28][2]  ( .D(datain[2]), .E(n1083), .CK(clk), .QN(n326) );
  EDFFX1 \data_reg[28][1]  ( .D(datain[1]), .E(n1083), .CK(clk), .QN(n327) );
  EDFFX1 \data_reg[28][0]  ( .D(datain[0]), .E(n1083), .CK(clk), .QN(n328) );
  EDFFX1 \data_reg[29][7]  ( .D(datain[7]), .E(n1084), .CK(clk), .QN(n329) );
  EDFFX1 \data_reg[29][6]  ( .D(datain[6]), .E(n1084), .CK(clk), .QN(n330) );
  EDFFX1 \data_reg[29][5]  ( .D(datain[5]), .E(n1084), .CK(clk), .QN(n331) );
  EDFFX1 \data_reg[29][4]  ( .D(datain[4]), .E(n1084), .CK(clk), .QN(n332) );
  EDFFX1 \data_reg[29][3]  ( .D(datain[3]), .E(n1084), .CK(clk), .QN(n333) );
  EDFFX1 \data_reg[29][2]  ( .D(datain[2]), .E(n1084), .CK(clk), .QN(n334) );
  EDFFX1 \data_reg[29][1]  ( .D(datain[1]), .E(n1084), .CK(clk), .QN(n335) );
  EDFFX1 \data_reg[29][0]  ( .D(datain[0]), .E(n1084), .CK(clk), .QN(n336) );
  EDFFX1 \data_reg[30][7]  ( .D(datain[7]), .E(n1085), .CK(clk), .QN(n337) );
  EDFFX1 \data_reg[30][6]  ( .D(datain[6]), .E(n1085), .CK(clk), .QN(n338) );
  EDFFX1 \data_reg[30][5]  ( .D(datain[5]), .E(n1085), .CK(clk), .QN(n339) );
  EDFFX1 \data_reg[30][4]  ( .D(datain[4]), .E(n1085), .CK(clk), .QN(n340) );
  EDFFX1 \data_reg[30][3]  ( .D(datain[3]), .E(n1085), .CK(clk), .QN(n341) );
  EDFFX1 \data_reg[30][2]  ( .D(datain[2]), .E(n1085), .CK(clk), .QN(n342) );
  EDFFX1 \data_reg[30][1]  ( .D(datain[1]), .E(n1085), .CK(clk), .QN(n343) );
  EDFFX1 \data_reg[30][0]  ( .D(datain[0]), .E(n1085), .CK(clk), .QN(n344) );
  EDFFX1 \data_reg[31][7]  ( .D(datain[7]), .E(n1086), .CK(clk), .QN(n345) );
  EDFFX1 \data_reg[31][6]  ( .D(datain[6]), .E(n1086), .CK(clk), .QN(n346) );
  EDFFX1 \data_reg[31][5]  ( .D(datain[5]), .E(n1086), .CK(clk), .QN(n347) );
  EDFFX1 \data_reg[31][4]  ( .D(datain[4]), .E(n1086), .CK(clk), .QN(n348) );
  EDFFX1 \data_reg[31][3]  ( .D(datain[3]), .E(n1086), .CK(clk), .QN(n349) );
  EDFFX1 \data_reg[31][2]  ( .D(datain[2]), .E(n1086), .CK(clk), .QN(n350) );
  EDFFX1 \data_reg[31][1]  ( .D(datain[1]), .E(n1086), .CK(clk), .QN(n351) );
  EDFFX1 \data_reg[31][0]  ( .D(datain[0]), .E(n1086), .CK(clk), .QN(n352) );
  EDFFX1 \data_reg[32][7]  ( .D(datain[7]), .E(n1087), .CK(clk), .QN(n353) );
  EDFFX1 \data_reg[32][6]  ( .D(datain[6]), .E(n1087), .CK(clk), .QN(n354) );
  EDFFX1 \data_reg[32][5]  ( .D(datain[5]), .E(n1087), .CK(clk), .QN(n355) );
  EDFFX1 \data_reg[32][4]  ( .D(datain[4]), .E(n1087), .CK(clk), .QN(n356) );
  EDFFX1 \data_reg[32][3]  ( .D(datain[3]), .E(n1087), .CK(clk), .QN(n357) );
  EDFFX1 \data_reg[32][2]  ( .D(datain[2]), .E(n1087), .CK(clk), .QN(n358) );
  EDFFX1 \data_reg[32][1]  ( .D(datain[1]), .E(n1087), .CK(clk), .QN(n359) );
  EDFFX1 \data_reg[32][0]  ( .D(datain[0]), .E(n1087), .CK(clk), .QN(n360) );
  EDFFX1 \data_reg[33][7]  ( .D(datain[7]), .E(n1088), .CK(clk), .QN(n361) );
  EDFFX1 \data_reg[33][6]  ( .D(datain[6]), .E(n1088), .CK(clk), .QN(n362) );
  EDFFX1 \data_reg[33][5]  ( .D(datain[5]), .E(n1088), .CK(clk), .QN(n363) );
  EDFFX1 \data_reg[33][4]  ( .D(datain[4]), .E(n1088), .CK(clk), .QN(n364) );
  EDFFX1 \data_reg[33][3]  ( .D(datain[3]), .E(n1088), .CK(clk), .QN(n365) );
  EDFFX1 \data_reg[33][2]  ( .D(datain[2]), .E(n1088), .CK(clk), .QN(n366) );
  EDFFX1 \data_reg[33][1]  ( .D(datain[1]), .E(n1088), .CK(clk), .QN(n367) );
  EDFFX1 \data_reg[33][0]  ( .D(datain[0]), .E(n1088), .CK(clk), .QN(n368) );
  EDFFX1 \data_reg[34][7]  ( .D(datain[7]), .E(n1089), .CK(clk), .QN(n369) );
  EDFFX1 \data_reg[34][6]  ( .D(datain[6]), .E(n1089), .CK(clk), .QN(n370) );
  EDFFX1 \data_reg[34][5]  ( .D(datain[5]), .E(n1089), .CK(clk), .QN(n371) );
  EDFFX1 \data_reg[34][4]  ( .D(datain[4]), .E(n1089), .CK(clk), .QN(n372) );
  EDFFX1 \data_reg[34][3]  ( .D(datain[3]), .E(n1089), .CK(clk), .QN(n373) );
  EDFFX1 \data_reg[34][2]  ( .D(datain[2]), .E(n1089), .CK(clk), .QN(n374) );
  EDFFX1 \data_reg[34][1]  ( .D(datain[1]), .E(n1089), .CK(clk), .QN(n375) );
  EDFFX1 \data_reg[34][0]  ( .D(datain[0]), .E(n1089), .CK(clk), .QN(n376) );
  EDFFX1 \data_reg[35][7]  ( .D(datain[7]), .E(n1090), .CK(clk), .QN(n377) );
  EDFFX1 \data_reg[35][6]  ( .D(datain[6]), .E(n1090), .CK(clk), .QN(n378) );
  EDFFX1 \data_reg[35][5]  ( .D(datain[5]), .E(n1090), .CK(clk), .QN(n379) );
  EDFFX1 \data_reg[35][4]  ( .D(datain[4]), .E(n1090), .CK(clk), .QN(n380) );
  EDFFX1 \data_reg[35][3]  ( .D(datain[3]), .E(n1090), .CK(clk), .QN(n381) );
  EDFFX1 \data_reg[35][2]  ( .D(datain[2]), .E(n1090), .CK(clk), .QN(n382) );
  EDFFX1 \data_reg[35][1]  ( .D(datain[1]), .E(n1090), .CK(clk), .QN(n383) );
  EDFFX1 \data_reg[35][0]  ( .D(datain[0]), .E(n1090), .CK(clk), .QN(n384) );
  DFFRXL \col_reg[0]  ( .D(n728), .CK(clk), .RN(n1054), .QN(n386) );
  DFFSXL \col_reg[1]  ( .D(n727), .CK(clk), .SN(n1054), .QN(n385) );
  DFFRXL output_valid_reg ( .D(n732), .CK(clk), .RN(n1054), .Q(output_valid), 
        .QN(n1053) );
  DFFRXL busy_reg ( .D(n731), .CK(clk), .RN(n1054), .Q(busy), .QN(n1052) );
  DFFSXL \row_reg[1]  ( .D(n729), .CK(clk), .SN(n1054), .Q(row[1]), .QN(n748)
         );
  DFFRXL \dataout_reg[0]  ( .D(n719), .CK(clk), .RN(n1054), .Q(dataout[0]) );
  DFFRXL \dataout_reg[1]  ( .D(n720), .CK(clk), .RN(n1054), .Q(dataout[1]) );
  DFFRXL \dataout_reg[2]  ( .D(n721), .CK(clk), .RN(n1054), .Q(dataout[2]) );
  DFFRXL \dataout_reg[3]  ( .D(n722), .CK(clk), .RN(n1054), .Q(dataout[3]) );
  DFFRXL \dataout_reg[4]  ( .D(n723), .CK(clk), .RN(n1054), .Q(dataout[4]) );
  DFFRXL \dataout_reg[5]  ( .D(n724), .CK(clk), .RN(n1054), .Q(dataout[5]) );
  DFFRXL \dataout_reg[6]  ( .D(n725), .CK(clk), .RN(n1054), .Q(dataout[6]) );
  DFFRXL \dataout_reg[7]  ( .D(n726), .CK(clk), .RN(n1054), .Q(dataout[7]) );
  DFFRXL \row_reg[0]  ( .D(n730), .CK(clk), .RN(n1054), .Q(row[0]), .QN(n746)
         );
  DFFRXL \cnt_reg[0]  ( .D(n741), .CK(clk), .RN(n1054), .Q(cnt[0]), .QN(n96)
         );
  DFFRXL \cnt_reg[4]  ( .D(n733), .CK(clk), .RN(n1054), .Q(cnt[4]), .QN(n92)
         );
  DFFRXL \cnt_reg[1]  ( .D(n736), .CK(clk), .RN(n1054), .Q(cnt[1]), .QN(n95)
         );
  DFFRXL \cnt_reg[2]  ( .D(n735), .CK(clk), .RN(n1054), .Q(cnt[2]), .QN(n94)
         );
  DFFRXL \cnt_reg[3]  ( .D(n734), .CK(clk), .RN(n1054), .Q(cnt[3]), .QN(n93)
         );
  ADDHXL \r407/U1_1_4  ( .A(cnt[4]), .B(\r407/carry[4] ), .CO(\r407/carry[5] ), 
        .S(N201) );
  ADDHXL \r407/U1_1_1  ( .A(cnt[1]), .B(cnt[0]), .CO(\r407/carry[2] ), .S(N198) );
  ADDHXL \r407/U1_1_3  ( .A(cnt[3]), .B(\r407/carry[3] ), .CO(\r407/carry[4] ), 
        .S(N200) );
  ADDHXL \r407/U1_1_2  ( .A(cnt[2]), .B(\r407/carry[2] ), .CO(\r407/carry[3] ), 
        .S(N199) );
  ADDFXL \add_0_root_add_171_2/U1_2  ( .A(\col_t[2] ), .B(N450), .CI(
        \add_0_root_add_171_2/carry[2] ), .CO(\add_0_root_add_171_2/carry[3] ), 
        .S(outpos[2]) );
  ADDFXL \add_1_root_add_171_2/U1_3  ( .A(row_t[1]), .B(row_t[2]), .CI(
        \add_1_root_add_171_2/carry[3] ), .CO(\add_1_root_add_171_2/carry[4] ), 
        .S(N451) );
  OR2X1 U414 ( .A(n752), .B(n753), .Y(n749) );
  INVX3 U415 ( .A(reset), .Y(n1054) );
  XNOR2X1 U416 ( .A(N452), .B(n749), .Y(outpos[4]) );
  XNOR2X1 U417 ( .A(n750), .B(\add_0_root_add_171_2/carry[5] ), .Y(outpos[5])
         );
  OR2X1 U418 ( .A(n757), .B(n758), .Y(n750) );
  NOR2X1 U419 ( .A(n754), .B(n749), .Y(\add_0_root_add_171_2/carry[5] ) );
  XNOR2X1 U420 ( .A(N451), .B(n753), .Y(outpos[3]) );
  CLKINVX1 U421 ( .A(N452), .Y(n754) );
  CLKINVX1 U422 ( .A(\add_1_root_add_171_2/carry[4] ), .Y(n757) );
  CLKINVX1 U423 ( .A(N451), .Y(n752) );
  XNOR2X1 U424 ( .A(row_t[2]), .B(n757), .Y(N452) );
  XNOR2X1 U425 ( .A(N449), .B(n751), .Y(outpos[1]) );
  CLKINVX1 U426 ( .A(N449), .Y(n755) );
  CLKINVX1 U427 ( .A(row_t[2]), .Y(n758) );
  NOR2X1 U428 ( .A(n755), .B(n756), .Y(\add_1_root_add_171_2/carry[3] ) );
  CLKINVX1 U429 ( .A(row_t[1]), .Y(n756) );
  CLKINVX1 U430 ( .A(\add_0_root_add_171_2/carry[3] ), .Y(n753) );
  XOR2X1 U431 ( .A(n1049), .B(n1051), .Y(n751) );
  NOR2X1 U432 ( .A(n755), .B(n751), .Y(\add_0_root_add_171_2/carry[2] ) );
  XNOR2X1 U433 ( .A(row_t[1]), .B(n755), .Y(N450) );
  XNOR2X1 U434 ( .A(n91), .B(n759), .Y(row_t[2]) );
  OAI21XL U435 ( .A0(n92), .A1(n760), .B0(n761), .Y(n759) );
  OAI21XL U436 ( .A0(n762), .A1(cnt[4]), .B0(row[1]), .Y(n761) );
  CLKINVX1 U437 ( .A(n762), .Y(n760) );
  XNOR2X1 U438 ( .A(n762), .B(n763), .Y(row_t[1]) );
  XNOR2X1 U439 ( .A(n748), .B(n92), .Y(n763) );
  NOR2X1 U440 ( .A(n746), .B(n93), .Y(n762) );
  OAI2BB1X1 U441 ( .A0N(n744), .A1N(n764), .B0(n765), .Y(next) );
  NOR2X1 U442 ( .A(n766), .B(n767), .Y(n1055) );
  NOR2X1 U443 ( .A(n766), .B(n768), .Y(n1056) );
  NOR2X1 U444 ( .A(n769), .B(n766), .Y(n1057) );
  NOR2X1 U445 ( .A(n766), .B(n770), .Y(n1058) );
  NOR2X1 U446 ( .A(n766), .B(n771), .Y(n1059) );
  NOR2X1 U447 ( .A(n766), .B(n772), .Y(n1060) );
  NOR2X1 U448 ( .A(n766), .B(n773), .Y(n1061) );
  NOR2X1 U449 ( .A(n766), .B(n774), .Y(n1062) );
  NAND2X1 U450 ( .A(n775), .B(n776), .Y(n766) );
  NOR2X1 U451 ( .A(n767), .B(n777), .Y(n1063) );
  NOR2X1 U452 ( .A(n768), .B(n777), .Y(n1064) );
  NOR2X1 U453 ( .A(n769), .B(n777), .Y(n1065) );
  NOR2X1 U454 ( .A(n770), .B(n777), .Y(n1066) );
  NOR2X1 U455 ( .A(n771), .B(n777), .Y(n1067) );
  NOR2X1 U456 ( .A(n772), .B(n777), .Y(n1068) );
  NOR2X1 U457 ( .A(n773), .B(n777), .Y(n1069) );
  NOR2X1 U458 ( .A(n774), .B(n777), .Y(n1070) );
  NAND3X1 U459 ( .A(n92), .B(cnt[3]), .C(n775), .Y(n777) );
  NOR2X1 U460 ( .A(n767), .B(n778), .Y(n1071) );
  NOR2X1 U461 ( .A(n768), .B(n778), .Y(n1072) );
  NOR2X1 U462 ( .A(n769), .B(n778), .Y(n1073) );
  NOR2X1 U463 ( .A(n770), .B(n778), .Y(n1074) );
  NOR2X1 U464 ( .A(n771), .B(n778), .Y(n1075) );
  NOR2X1 U465 ( .A(n772), .B(n778), .Y(n1076) );
  NOR2X1 U466 ( .A(n773), .B(n778), .Y(n1077) );
  NOR2X1 U467 ( .A(n774), .B(n778), .Y(n1078) );
  NAND3X1 U468 ( .A(n93), .B(cnt[4]), .C(n775), .Y(n778) );
  NOR2X1 U469 ( .A(n767), .B(n779), .Y(n1079) );
  NOR2X1 U470 ( .A(n768), .B(n779), .Y(n1080) );
  NOR2X1 U471 ( .A(n769), .B(n779), .Y(n1081) );
  NOR2X1 U472 ( .A(n770), .B(n779), .Y(n1082) );
  NOR2X1 U473 ( .A(n771), .B(n779), .Y(n1083) );
  NAND3X1 U474 ( .A(n96), .B(cnt[2]), .C(n95), .Y(n771) );
  NOR2X1 U475 ( .A(n772), .B(n779), .Y(n1084) );
  NAND3X1 U476 ( .A(cnt[2]), .B(cnt[0]), .C(n95), .Y(n772) );
  NOR2X1 U477 ( .A(n773), .B(n779), .Y(n1085) );
  NAND3X1 U478 ( .A(cnt[2]), .B(cnt[1]), .C(n96), .Y(n773) );
  NOR2X1 U479 ( .A(n774), .B(n779), .Y(n1086) );
  NAND3X1 U480 ( .A(cnt[4]), .B(cnt[3]), .C(n775), .Y(n779) );
  NOR2X1 U481 ( .A(n780), .B(n745), .Y(n775) );
  NAND3X1 U482 ( .A(cnt[1]), .B(cnt[0]), .C(cnt[2]), .Y(n774) );
  NOR2X1 U483 ( .A(n767), .B(n781), .Y(n1087) );
  NAND3X1 U484 ( .A(n96), .B(n94), .C(n95), .Y(n767) );
  NOR2X1 U485 ( .A(n768), .B(n781), .Y(n1088) );
  NAND3X1 U486 ( .A(n94), .B(cnt[0]), .C(n95), .Y(n768) );
  NOR2X1 U487 ( .A(n769), .B(n781), .Y(n1089) );
  NAND3BX1 U488 ( .AN(n780), .B(n745), .C(n776), .Y(n781) );
  NOR2X1 U489 ( .A(n780), .B(n782), .Y(n1090) );
  NAND2X1 U490 ( .A(n783), .B(n1054), .Y(n780) );
  MXI2X1 U491 ( .A(n784), .B(n785), .S0(cnt[0]), .Y(n741) );
  MXI2X1 U492 ( .A(n786), .B(n787), .S0(n745), .Y(n740) );
  AOI221XL U493 ( .A0(n788), .A1(n92), .B0(n789), .B1(n790), .C0(n791), .Y(
        n787) );
  CLKINVX1 U494 ( .A(\r407/carry[5] ), .Y(n790) );
  AOI32X1 U495 ( .A0(cnt[4]), .A1(cnt[3]), .A2(n788), .B0(\r407/carry[5] ), 
        .B1(n789), .Y(n786) );
  OAI2BB2XL U496 ( .B0(n84), .B1(n792), .A0N(cmd[2]), .A1N(n793), .Y(n739) );
  OAI2BB2XL U497 ( .B0(n86), .B1(n792), .A0N(cmd[0]), .A1N(n793), .Y(n738) );
  OAI2BB2XL U498 ( .B0(n85), .B1(n792), .A0N(cmd[1]), .A1N(n793), .Y(n737) );
  AND2X1 U499 ( .A(n792), .B(n78), .Y(n793) );
  OAI211X1 U500 ( .A0(n794), .A1(n782), .B0(n795), .C0(n765), .Y(n792) );
  AO21X1 U501 ( .A0(n796), .A1(n797), .B0(n78), .Y(n795) );
  OAI2BB2XL U502 ( .B0(n785), .B1(n95), .A0N(N198), .A1N(n789), .Y(n736) );
  OAI2BB2XL U503 ( .B0(n785), .B1(n94), .A0N(N199), .A1N(n789), .Y(n735) );
  OAI211X1 U504 ( .A0(n93), .A1(n785), .B0(n798), .C0(n799), .Y(n734) );
  NAND2X1 U505 ( .A(N200), .B(n789), .Y(n799) );
  OAI2BB1X1 U506 ( .A0N(N201), .A1N(n789), .B0(n800), .Y(n733) );
  MXI2X1 U507 ( .A(n801), .B(n791), .S0(cnt[4]), .Y(n800) );
  NAND2X1 U508 ( .A(n785), .B(n798), .Y(n791) );
  NAND2X1 U509 ( .A(n788), .B(n93), .Y(n798) );
  NAND3BX1 U510 ( .AN(n802), .B(n744), .C(n803), .Y(n785) );
  AND2X1 U511 ( .A(n788), .B(cnt[3]), .Y(n801) );
  NOR2X1 U512 ( .A(n804), .B(n769), .Y(n788) );
  CLKINVX1 U513 ( .A(n784), .Y(n789) );
  AOI22X1 U514 ( .A0(n769), .A1(n805), .B0(n782), .B1(n783), .Y(n784) );
  NAND3BX1 U515 ( .AN(n770), .B(n776), .C(n745), .Y(n782) );
  NOR2X1 U516 ( .A(cnt[3]), .B(cnt[4]), .Y(n776) );
  NAND3X1 U517 ( .A(cnt[1]), .B(cnt[0]), .C(n94), .Y(n770) );
  CLKINVX1 U518 ( .A(n804), .Y(n805) );
  OAI21XL U519 ( .A0(n78), .A1(n1053), .B0(n804), .Y(n732) );
  OAI21XL U520 ( .A0(n1052), .A1(n806), .B0(n765), .Y(n731) );
  NAND2X1 U521 ( .A(n78), .B(cmd_valid), .Y(n765) );
  NOR2X1 U522 ( .A(n764), .B(n78), .Y(n806) );
  NAND3X1 U523 ( .A(n93), .B(n802), .C(n807), .Y(n764) );
  NOR3X1 U524 ( .A(n769), .B(n92), .C(n745), .Y(n807) );
  NAND3X1 U525 ( .A(n94), .B(cnt[1]), .C(n96), .Y(n769) );
  MXI2X1 U526 ( .A(n808), .B(n809), .S0(n746), .Y(n730) );
  OAI21XL U527 ( .A0(n810), .A1(n811), .B0(n812), .Y(n809) );
  OA21XL U528 ( .A0(n813), .A1(n814), .B0(n812), .Y(n808) );
  OAI22XL U529 ( .A0(n815), .A1(n816), .B0(n817), .B1(n748), .Y(n729) );
  NOR3X1 U530 ( .A(row[0]), .B(n810), .C(n815), .Y(n817) );
  OA21XL U531 ( .A0(n746), .A1(n811), .B0(n803), .Y(n816) );
  CLKINVX1 U532 ( .A(n812), .Y(n815) );
  OAI21XL U533 ( .A0(n797), .A1(n78), .B0(n794), .Y(n812) );
  MXI2X1 U534 ( .A(n818), .B(n819), .S0(n386), .Y(n728) );
  OAI21XL U535 ( .A0(n820), .A1(n811), .B0(n821), .Y(n819) );
  OA21XL U536 ( .A0(n813), .A1(n822), .B0(n821), .Y(n818) );
  CLKINVX1 U537 ( .A(n811), .Y(n813) );
  OAI22XL U538 ( .A0(n823), .A1(n824), .B0(n385), .B1(n825), .Y(n727) );
  NOR3BXL U539 ( .AN(n386), .B(n820), .C(n823), .Y(n825) );
  OA21XL U540 ( .A0(n811), .A1(n386), .B0(n803), .Y(n824) );
  OAI221XL U541 ( .A0(n797), .A1(n748), .B0(n385), .B1(n796), .C0(n826), .Y(
        n811) );
  NAND3X1 U542 ( .A(n814), .B(n822), .C(n827), .Y(n826) );
  OAI22XL U543 ( .A0(n386), .A1(n796), .B0(n797), .B1(n746), .Y(n827) );
  CLKINVX1 U544 ( .A(n820), .Y(n822) );
  NOR2X1 U545 ( .A(n743), .B(n742), .Y(n820) );
  CLKINVX1 U546 ( .A(n810), .Y(n814) );
  NOR2X1 U547 ( .A(n84), .B(n86), .Y(n810) );
  NAND2X1 U548 ( .A(n85), .B(n742), .Y(n797) );
  CLKINVX1 U549 ( .A(n821), .Y(n823) );
  OAI21XL U550 ( .A0(n796), .A1(n78), .B0(n794), .Y(n821) );
  CLKINVX1 U551 ( .A(n783), .Y(n794) );
  NOR2X1 U552 ( .A(n803), .B(n78), .Y(n783) );
  NAND3X1 U553 ( .A(n84), .B(n743), .C(n85), .Y(n803) );
  NAND2X1 U554 ( .A(n84), .B(n747), .Y(n796) );
  CLKMX2X2 U555 ( .A(n828), .B(dataout[7]), .S0(n804), .Y(n726) );
  NAND4X1 U556 ( .A(n829), .B(n830), .C(n831), .D(n832), .Y(n828) );
  NOR4X1 U557 ( .A(n833), .B(n834), .C(n835), .D(n836), .Y(n832) );
  OAI22XL U558 ( .A0(n837), .A1(n369), .B0(n838), .B1(n377), .Y(n836) );
  OAI22XL U559 ( .A0(n839), .A1(n361), .B0(n840), .B1(n345), .Y(n835) );
  OAI22XL U560 ( .A0(n841), .A1(n353), .B0(n842), .B1(n329), .Y(n834) );
  OAI222XL U561 ( .A0(n843), .A1(n313), .B0(n844), .B1(n321), .C0(n845), .C1(
        n337), .Y(n833) );
  NOR4X1 U562 ( .A(n846), .B(n847), .C(n848), .D(n849), .Y(n831) );
  OAI22XL U563 ( .A0(n850), .A1(n297), .B0(n851), .B1(n305), .Y(n849) );
  OAI22XL U564 ( .A0(n852), .A1(n289), .B0(n853), .B1(n273), .Y(n848) );
  OAI22XL U565 ( .A0(n854), .A1(n281), .B0(n855), .B1(n257), .Y(n847) );
  OAI222XL U566 ( .A0(n856), .A1(n241), .B0(n857), .B1(n249), .C0(n858), .C1(
        n265), .Y(n846) );
  NOR4X1 U567 ( .A(n859), .B(n860), .C(n861), .D(n862), .Y(n830) );
  OAI22XL U568 ( .A0(n863), .A1(n225), .B0(n864), .B1(n233), .Y(n862) );
  OAI22XL U569 ( .A0(n865), .A1(n217), .B0(n866), .B1(n201), .Y(n861) );
  OAI22XL U570 ( .A0(n867), .A1(n209), .B0(n868), .B1(n185), .Y(n860) );
  OAI222XL U571 ( .A0(n869), .A1(n169), .B0(n870), .B1(n177), .C0(n871), .C1(
        n193), .Y(n859) );
  NOR4X1 U572 ( .A(n872), .B(n873), .C(n874), .D(n875), .Y(n829) );
  OAI22XL U573 ( .A0(n876), .A1(n153), .B0(n877), .B1(n161), .Y(n875) );
  OAI22XL U574 ( .A0(n878), .A1(n145), .B0(n879), .B1(n129), .Y(n874) );
  OAI22XL U575 ( .A0(n880), .A1(n137), .B0(n881), .B1(n113), .Y(n873) );
  OAI222XL U576 ( .A0(n882), .A1(n97), .B0(n883), .B1(n105), .C0(n884), .C1(
        n121), .Y(n872) );
  CLKMX2X2 U577 ( .A(n885), .B(dataout[6]), .S0(n804), .Y(n725) );
  NAND4X1 U578 ( .A(n886), .B(n887), .C(n888), .D(n889), .Y(n885) );
  NOR4X1 U579 ( .A(n890), .B(n891), .C(n892), .D(n893), .Y(n889) );
  OAI22XL U580 ( .A0(n837), .A1(n370), .B0(n838), .B1(n378), .Y(n893) );
  OAI22XL U581 ( .A0(n839), .A1(n362), .B0(n840), .B1(n346), .Y(n892) );
  OAI22XL U582 ( .A0(n841), .A1(n354), .B0(n842), .B1(n330), .Y(n891) );
  OAI222XL U583 ( .A0(n843), .A1(n314), .B0(n844), .B1(n322), .C0(n845), .C1(
        n338), .Y(n890) );
  NOR4X1 U584 ( .A(n894), .B(n895), .C(n896), .D(n897), .Y(n888) );
  OAI22XL U585 ( .A0(n850), .A1(n298), .B0(n851), .B1(n306), .Y(n897) );
  OAI22XL U586 ( .A0(n852), .A1(n290), .B0(n853), .B1(n274), .Y(n896) );
  OAI22XL U587 ( .A0(n854), .A1(n282), .B0(n855), .B1(n258), .Y(n895) );
  OAI222XL U588 ( .A0(n856), .A1(n242), .B0(n857), .B1(n250), .C0(n858), .C1(
        n266), .Y(n894) );
  NOR4X1 U589 ( .A(n898), .B(n899), .C(n900), .D(n901), .Y(n887) );
  OAI22XL U590 ( .A0(n863), .A1(n226), .B0(n864), .B1(n234), .Y(n901) );
  OAI22XL U591 ( .A0(n865), .A1(n218), .B0(n866), .B1(n202), .Y(n900) );
  OAI22XL U592 ( .A0(n867), .A1(n210), .B0(n868), .B1(n186), .Y(n899) );
  OAI222XL U593 ( .A0(n869), .A1(n170), .B0(n870), .B1(n178), .C0(n871), .C1(
        n194), .Y(n898) );
  NOR4X1 U594 ( .A(n902), .B(n903), .C(n904), .D(n905), .Y(n886) );
  OAI22XL U595 ( .A0(n876), .A1(n154), .B0(n877), .B1(n162), .Y(n905) );
  OAI22XL U596 ( .A0(n878), .A1(n146), .B0(n879), .B1(n130), .Y(n904) );
  OAI22XL U597 ( .A0(n880), .A1(n138), .B0(n881), .B1(n114), .Y(n903) );
  OAI222XL U598 ( .A0(n882), .A1(n98), .B0(n883), .B1(n106), .C0(n884), .C1(
        n122), .Y(n902) );
  CLKMX2X2 U599 ( .A(n906), .B(dataout[5]), .S0(n804), .Y(n724) );
  NAND4X1 U600 ( .A(n907), .B(n908), .C(n909), .D(n910), .Y(n906) );
  NOR4X1 U601 ( .A(n911), .B(n912), .C(n913), .D(n914), .Y(n910) );
  OAI22XL U602 ( .A0(n837), .A1(n371), .B0(n838), .B1(n379), .Y(n914) );
  OAI22XL U603 ( .A0(n839), .A1(n363), .B0(n840), .B1(n347), .Y(n913) );
  OAI22XL U604 ( .A0(n841), .A1(n355), .B0(n842), .B1(n331), .Y(n912) );
  OAI222XL U605 ( .A0(n843), .A1(n315), .B0(n844), .B1(n323), .C0(n845), .C1(
        n339), .Y(n911) );
  NOR4X1 U606 ( .A(n915), .B(n916), .C(n917), .D(n918), .Y(n909) );
  OAI22XL U607 ( .A0(n850), .A1(n299), .B0(n851), .B1(n307), .Y(n918) );
  OAI22XL U608 ( .A0(n852), .A1(n291), .B0(n853), .B1(n275), .Y(n917) );
  OAI22XL U609 ( .A0(n854), .A1(n283), .B0(n855), .B1(n259), .Y(n916) );
  OAI222XL U610 ( .A0(n856), .A1(n243), .B0(n857), .B1(n251), .C0(n858), .C1(
        n267), .Y(n915) );
  NOR4X1 U611 ( .A(n919), .B(n920), .C(n921), .D(n922), .Y(n908) );
  OAI22XL U612 ( .A0(n863), .A1(n227), .B0(n864), .B1(n235), .Y(n922) );
  OAI22XL U613 ( .A0(n865), .A1(n219), .B0(n866), .B1(n203), .Y(n921) );
  OAI22XL U614 ( .A0(n867), .A1(n211), .B0(n868), .B1(n187), .Y(n920) );
  OAI222XL U615 ( .A0(n869), .A1(n171), .B0(n870), .B1(n179), .C0(n871), .C1(
        n195), .Y(n919) );
  NOR4X1 U616 ( .A(n923), .B(n924), .C(n925), .D(n926), .Y(n907) );
  OAI22XL U617 ( .A0(n876), .A1(n155), .B0(n877), .B1(n163), .Y(n926) );
  OAI22XL U618 ( .A0(n878), .A1(n147), .B0(n879), .B1(n131), .Y(n925) );
  OAI22XL U619 ( .A0(n880), .A1(n139), .B0(n881), .B1(n115), .Y(n924) );
  OAI222XL U620 ( .A0(n882), .A1(n99), .B0(n883), .B1(n107), .C0(n884), .C1(
        n123), .Y(n923) );
  CLKMX2X2 U621 ( .A(n927), .B(dataout[4]), .S0(n804), .Y(n723) );
  NAND4X1 U622 ( .A(n928), .B(n929), .C(n930), .D(n931), .Y(n927) );
  NOR4X1 U623 ( .A(n932), .B(n933), .C(n934), .D(n935), .Y(n931) );
  OAI22XL U624 ( .A0(n837), .A1(n372), .B0(n838), .B1(n380), .Y(n935) );
  OAI22XL U625 ( .A0(n839), .A1(n364), .B0(n840), .B1(n348), .Y(n934) );
  OAI22XL U626 ( .A0(n841), .A1(n356), .B0(n842), .B1(n332), .Y(n933) );
  OAI222XL U627 ( .A0(n843), .A1(n316), .B0(n844), .B1(n324), .C0(n845), .C1(
        n340), .Y(n932) );
  NOR4X1 U628 ( .A(n936), .B(n937), .C(n938), .D(n939), .Y(n930) );
  OAI22XL U629 ( .A0(n850), .A1(n300), .B0(n851), .B1(n308), .Y(n939) );
  OAI22XL U630 ( .A0(n852), .A1(n292), .B0(n853), .B1(n276), .Y(n938) );
  OAI22XL U631 ( .A0(n854), .A1(n284), .B0(n855), .B1(n260), .Y(n937) );
  OAI222XL U632 ( .A0(n856), .A1(n244), .B0(n857), .B1(n252), .C0(n858), .C1(
        n268), .Y(n936) );
  NOR4X1 U633 ( .A(n940), .B(n941), .C(n942), .D(n943), .Y(n929) );
  OAI22XL U634 ( .A0(n863), .A1(n228), .B0(n864), .B1(n236), .Y(n943) );
  OAI22XL U635 ( .A0(n865), .A1(n220), .B0(n866), .B1(n204), .Y(n942) );
  OAI22XL U636 ( .A0(n867), .A1(n212), .B0(n868), .B1(n188), .Y(n941) );
  OAI222XL U637 ( .A0(n869), .A1(n172), .B0(n870), .B1(n180), .C0(n871), .C1(
        n196), .Y(n940) );
  NOR4X1 U638 ( .A(n944), .B(n945), .C(n946), .D(n947), .Y(n928) );
  OAI22XL U639 ( .A0(n876), .A1(n156), .B0(n877), .B1(n164), .Y(n947) );
  OAI22XL U640 ( .A0(n878), .A1(n148), .B0(n879), .B1(n132), .Y(n946) );
  OAI22XL U641 ( .A0(n880), .A1(n140), .B0(n881), .B1(n116), .Y(n945) );
  OAI222XL U642 ( .A0(n882), .A1(n100), .B0(n883), .B1(n108), .C0(n884), .C1(
        n124), .Y(n944) );
  CLKMX2X2 U643 ( .A(n948), .B(dataout[3]), .S0(n804), .Y(n722) );
  NAND4X1 U644 ( .A(n949), .B(n950), .C(n951), .D(n952), .Y(n948) );
  NOR4X1 U645 ( .A(n953), .B(n954), .C(n955), .D(n956), .Y(n952) );
  OAI22XL U646 ( .A0(n837), .A1(n373), .B0(n838), .B1(n381), .Y(n956) );
  OAI22XL U647 ( .A0(n839), .A1(n365), .B0(n840), .B1(n349), .Y(n955) );
  OAI22XL U648 ( .A0(n841), .A1(n357), .B0(n842), .B1(n333), .Y(n954) );
  OAI222XL U649 ( .A0(n843), .A1(n317), .B0(n844), .B1(n325), .C0(n845), .C1(
        n341), .Y(n953) );
  NOR4X1 U650 ( .A(n957), .B(n958), .C(n959), .D(n960), .Y(n951) );
  OAI22XL U651 ( .A0(n850), .A1(n301), .B0(n851), .B1(n309), .Y(n960) );
  OAI22XL U652 ( .A0(n852), .A1(n293), .B0(n853), .B1(n277), .Y(n959) );
  OAI22XL U653 ( .A0(n854), .A1(n285), .B0(n855), .B1(n261), .Y(n958) );
  OAI222XL U654 ( .A0(n856), .A1(n245), .B0(n857), .B1(n253), .C0(n858), .C1(
        n269), .Y(n957) );
  NOR4X1 U655 ( .A(n961), .B(n962), .C(n963), .D(n964), .Y(n950) );
  OAI22XL U656 ( .A0(n863), .A1(n229), .B0(n864), .B1(n237), .Y(n964) );
  OAI22XL U657 ( .A0(n865), .A1(n221), .B0(n866), .B1(n205), .Y(n963) );
  OAI22XL U658 ( .A0(n867), .A1(n213), .B0(n868), .B1(n189), .Y(n962) );
  OAI222XL U659 ( .A0(n869), .A1(n173), .B0(n870), .B1(n181), .C0(n871), .C1(
        n197), .Y(n961) );
  NOR4X1 U660 ( .A(n965), .B(n966), .C(n967), .D(n968), .Y(n949) );
  OAI22XL U661 ( .A0(n876), .A1(n157), .B0(n877), .B1(n165), .Y(n968) );
  OAI22XL U662 ( .A0(n878), .A1(n149), .B0(n879), .B1(n133), .Y(n967) );
  OAI22XL U663 ( .A0(n880), .A1(n141), .B0(n881), .B1(n117), .Y(n966) );
  OAI222XL U664 ( .A0(n882), .A1(n101), .B0(n883), .B1(n109), .C0(n884), .C1(
        n125), .Y(n965) );
  CLKMX2X2 U665 ( .A(n969), .B(dataout[2]), .S0(n804), .Y(n721) );
  NAND4X1 U666 ( .A(n970), .B(n971), .C(n972), .D(n973), .Y(n969) );
  NOR4X1 U667 ( .A(n974), .B(n975), .C(n976), .D(n977), .Y(n973) );
  OAI22XL U668 ( .A0(n837), .A1(n374), .B0(n838), .B1(n382), .Y(n977) );
  OAI22XL U669 ( .A0(n839), .A1(n366), .B0(n840), .B1(n350), .Y(n976) );
  OAI22XL U670 ( .A0(n841), .A1(n358), .B0(n842), .B1(n334), .Y(n975) );
  OAI222XL U671 ( .A0(n843), .A1(n318), .B0(n844), .B1(n326), .C0(n845), .C1(
        n342), .Y(n974) );
  NOR4X1 U672 ( .A(n978), .B(n979), .C(n980), .D(n981), .Y(n972) );
  OAI22XL U673 ( .A0(n850), .A1(n302), .B0(n851), .B1(n310), .Y(n981) );
  OAI22XL U674 ( .A0(n852), .A1(n294), .B0(n853), .B1(n278), .Y(n980) );
  OAI22XL U675 ( .A0(n854), .A1(n286), .B0(n855), .B1(n262), .Y(n979) );
  OAI222XL U676 ( .A0(n856), .A1(n246), .B0(n857), .B1(n254), .C0(n858), .C1(
        n270), .Y(n978) );
  NOR4X1 U677 ( .A(n982), .B(n983), .C(n984), .D(n985), .Y(n971) );
  OAI22XL U678 ( .A0(n863), .A1(n230), .B0(n864), .B1(n238), .Y(n985) );
  OAI22XL U679 ( .A0(n865), .A1(n222), .B0(n866), .B1(n206), .Y(n984) );
  OAI22XL U680 ( .A0(n867), .A1(n214), .B0(n868), .B1(n190), .Y(n983) );
  OAI222XL U681 ( .A0(n869), .A1(n174), .B0(n870), .B1(n182), .C0(n871), .C1(
        n198), .Y(n982) );
  NOR4X1 U682 ( .A(n986), .B(n987), .C(n988), .D(n989), .Y(n970) );
  OAI22XL U683 ( .A0(n876), .A1(n158), .B0(n877), .B1(n166), .Y(n989) );
  OAI22XL U684 ( .A0(n878), .A1(n150), .B0(n879), .B1(n134), .Y(n988) );
  OAI22XL U685 ( .A0(n880), .A1(n142), .B0(n881), .B1(n118), .Y(n987) );
  OAI222XL U686 ( .A0(n882), .A1(n102), .B0(n883), .B1(n110), .C0(n884), .C1(
        n126), .Y(n986) );
  CLKMX2X2 U687 ( .A(n990), .B(dataout[1]), .S0(n804), .Y(n720) );
  NAND4X1 U688 ( .A(n991), .B(n992), .C(n993), .D(n994), .Y(n990) );
  NOR4X1 U689 ( .A(n995), .B(n996), .C(n997), .D(n998), .Y(n994) );
  OAI22XL U690 ( .A0(n837), .A1(n375), .B0(n838), .B1(n383), .Y(n998) );
  OAI22XL U691 ( .A0(n839), .A1(n367), .B0(n840), .B1(n351), .Y(n997) );
  OAI22XL U692 ( .A0(n841), .A1(n359), .B0(n842), .B1(n335), .Y(n996) );
  OAI222XL U693 ( .A0(n843), .A1(n319), .B0(n844), .B1(n327), .C0(n845), .C1(
        n343), .Y(n995) );
  NOR4X1 U694 ( .A(n999), .B(n1000), .C(n1001), .D(n1002), .Y(n993) );
  OAI22XL U695 ( .A0(n850), .A1(n303), .B0(n851), .B1(n311), .Y(n1002) );
  OAI22XL U696 ( .A0(n852), .A1(n295), .B0(n853), .B1(n279), .Y(n1001) );
  OAI22XL U697 ( .A0(n854), .A1(n287), .B0(n855), .B1(n263), .Y(n1000) );
  OAI222XL U698 ( .A0(n856), .A1(n247), .B0(n857), .B1(n255), .C0(n858), .C1(
        n271), .Y(n999) );
  NOR4X1 U699 ( .A(n1003), .B(n1004), .C(n1005), .D(n1006), .Y(n992) );
  OAI22XL U700 ( .A0(n863), .A1(n231), .B0(n864), .B1(n239), .Y(n1006) );
  OAI22XL U701 ( .A0(n865), .A1(n223), .B0(n866), .B1(n207), .Y(n1005) );
  OAI22XL U702 ( .A0(n867), .A1(n215), .B0(n868), .B1(n191), .Y(n1004) );
  OAI222XL U703 ( .A0(n869), .A1(n175), .B0(n870), .B1(n183), .C0(n871), .C1(
        n199), .Y(n1003) );
  NOR4X1 U704 ( .A(n1007), .B(n1008), .C(n1009), .D(n1010), .Y(n991) );
  OAI22XL U705 ( .A0(n876), .A1(n159), .B0(n877), .B1(n167), .Y(n1010) );
  OAI22XL U706 ( .A0(n878), .A1(n151), .B0(n879), .B1(n135), .Y(n1009) );
  OAI22XL U707 ( .A0(n880), .A1(n143), .B0(n881), .B1(n119), .Y(n1008) );
  OAI222XL U708 ( .A0(n882), .A1(n103), .B0(n883), .B1(n111), .C0(n884), .C1(
        n127), .Y(n1007) );
  CLKMX2X2 U709 ( .A(n1011), .B(dataout[0]), .S0(n804), .Y(n719) );
  NAND2X1 U710 ( .A(n802), .B(n744), .Y(n804) );
  NOR3X1 U711 ( .A(n747), .B(n742), .C(n743), .Y(n802) );
  NAND4X1 U712 ( .A(n1012), .B(n1013), .C(n1014), .D(n1015), .Y(n1011) );
  NOR4X1 U713 ( .A(n1016), .B(n1017), .C(n1018), .D(n1019), .Y(n1015) );
  OAI22XL U714 ( .A0(n837), .A1(n376), .B0(n838), .B1(n384), .Y(n1019) );
  NAND2X1 U715 ( .A(outpos[5]), .B(n1020), .Y(n838) );
  NAND2X1 U716 ( .A(outpos[5]), .B(n1021), .Y(n837) );
  OAI22XL U717 ( .A0(n839), .A1(n368), .B0(n840), .B1(n352), .Y(n1018) );
  NAND2X1 U718 ( .A(n1020), .B(n1022), .Y(n840) );
  NAND2X1 U719 ( .A(outpos[5]), .B(n1023), .Y(n839) );
  OAI22XL U720 ( .A0(n841), .A1(n360), .B0(n842), .B1(n336), .Y(n1017) );
  NAND2X1 U721 ( .A(n1023), .B(n1022), .Y(n842) );
  NAND2X1 U722 ( .A(outpos[5]), .B(n1024), .Y(n841) );
  OAI222XL U723 ( .A0(n843), .A1(n320), .B0(n844), .B1(n328), .C0(n845), .C1(
        n344), .Y(n1016) );
  NAND2X1 U724 ( .A(n1021), .B(n1022), .Y(n845) );
  NAND2X1 U725 ( .A(n1024), .B(n1022), .Y(n844) );
  AND3X1 U726 ( .A(outpos[4]), .B(outpos[3]), .C(outpos[2]), .Y(n1022) );
  NAND2X1 U727 ( .A(n1020), .B(n1025), .Y(n843) );
  NOR4X1 U728 ( .A(n1026), .B(n1027), .C(n1028), .D(n1029), .Y(n1014) );
  OAI22XL U729 ( .A0(n850), .A1(n304), .B0(n851), .B1(n312), .Y(n1029) );
  NAND2X1 U730 ( .A(n1021), .B(n1025), .Y(n851) );
  NAND2X1 U731 ( .A(n1023), .B(n1025), .Y(n850) );
  OAI22XL U732 ( .A0(n852), .A1(n296), .B0(n853), .B1(n280), .Y(n1028) );
  NAND2X1 U733 ( .A(n1030), .B(n1021), .Y(n853) );
  NAND2X1 U734 ( .A(n1025), .B(n1024), .Y(n852) );
  AND3X1 U735 ( .A(outpos[4]), .B(outpos[3]), .C(n1031), .Y(n1025) );
  OAI22XL U736 ( .A0(n854), .A1(n288), .B0(n855), .B1(n264), .Y(n1027) );
  NAND2X1 U737 ( .A(n1030), .B(n1024), .Y(n855) );
  NAND2X1 U738 ( .A(n1030), .B(n1020), .Y(n854) );
  OAI222XL U739 ( .A0(n856), .A1(n248), .B0(n857), .B1(n256), .C0(n858), .C1(
        n272), .Y(n1026) );
  NAND2X1 U740 ( .A(n1030), .B(n1023), .Y(n858) );
  AND3X1 U741 ( .A(outpos[4]), .B(outpos[2]), .C(n1032), .Y(n1030) );
  NAND2X1 U742 ( .A(n1033), .B(n1020), .Y(n857) );
  NAND2X1 U743 ( .A(n1033), .B(n1021), .Y(n856) );
  NOR4X1 U744 ( .A(n1034), .B(n1035), .C(n1036), .D(n1037), .Y(n1013) );
  OAI22XL U745 ( .A0(n863), .A1(n232), .B0(n864), .B1(n240), .Y(n1037) );
  NAND2X1 U746 ( .A(n1033), .B(n1023), .Y(n864) );
  NAND2X1 U747 ( .A(n1033), .B(n1024), .Y(n863) );
  AND3X1 U748 ( .A(outpos[4]), .B(n1031), .C(n1032), .Y(n1033) );
  OAI22XL U749 ( .A0(n865), .A1(n224), .B0(n866), .B1(n208), .Y(n1036) );
  NAND2X1 U750 ( .A(n1038), .B(n1023), .Y(n866) );
  NAND2X1 U751 ( .A(n1038), .B(n1020), .Y(n865) );
  OAI22XL U752 ( .A0(n867), .A1(n216), .B0(n868), .B1(n192), .Y(n1035) );
  NAND2X1 U753 ( .A(n1039), .B(n1020), .Y(n868) );
  NAND2X1 U754 ( .A(n1038), .B(n1021), .Y(n867) );
  OAI222XL U755 ( .A0(n869), .A1(n176), .B0(n870), .B1(n184), .C0(n871), .C1(
        n200), .Y(n1034) );
  NAND2X1 U756 ( .A(n1038), .B(n1024), .Y(n871) );
  NOR3X1 U757 ( .A(n1031), .B(outpos[4]), .C(n1032), .Y(n1038) );
  NAND2X1 U758 ( .A(n1039), .B(n1021), .Y(n870) );
  NAND2X1 U759 ( .A(n1039), .B(n1023), .Y(n869) );
  NOR4X1 U760 ( .A(n1040), .B(n1041), .C(n1042), .D(n1043), .Y(n1012) );
  OAI22XL U761 ( .A0(n876), .A1(n160), .B0(n877), .B1(n168), .Y(n1043) );
  NAND2X1 U762 ( .A(n1039), .B(n1024), .Y(n877) );
  NOR3X1 U763 ( .A(outpos[2]), .B(outpos[4]), .C(n1032), .Y(n1039) );
  CLKINVX1 U764 ( .A(outpos[3]), .Y(n1032) );
  NAND2X1 U765 ( .A(n1044), .B(n1020), .Y(n876) );
  OAI22XL U766 ( .A0(n878), .A1(n152), .B0(n879), .B1(n136), .Y(n1042) );
  NAND2X1 U767 ( .A(n1044), .B(n1024), .Y(n879) );
  NAND2X1 U768 ( .A(n1044), .B(n1021), .Y(n878) );
  OAI22XL U769 ( .A0(n880), .A1(n144), .B0(n881), .B1(n120), .Y(n1041) );
  NAND2X1 U770 ( .A(n1045), .B(n1021), .Y(n881) );
  AND2X1 U771 ( .A(outpos[1]), .B(n1046), .Y(n1021) );
  NAND2X1 U772 ( .A(n1044), .B(n1023), .Y(n880) );
  NOR3X1 U773 ( .A(outpos[3]), .B(outpos[4]), .C(n1031), .Y(n1044) );
  CLKINVX1 U774 ( .A(outpos[2]), .Y(n1031) );
  OAI222XL U775 ( .A0(n882), .A1(n104), .B0(n883), .B1(n112), .C0(n884), .C1(
        n128), .Y(n1040) );
  NAND2X1 U776 ( .A(n1045), .B(n1020), .Y(n884) );
  AND2X1 U777 ( .A(outpos[1]), .B(n1047), .Y(n1020) );
  NAND2X1 U778 ( .A(n1045), .B(n1023), .Y(n883) );
  NOR2X1 U779 ( .A(n1046), .B(outpos[1]), .Y(n1023) );
  NAND2X1 U780 ( .A(n1045), .B(n1024), .Y(n882) );
  NOR2X1 U781 ( .A(n1047), .B(outpos[1]), .Y(n1024) );
  CLKINVX1 U782 ( .A(n1046), .Y(n1047) );
  XOR2X1 U783 ( .A(n386), .B(cnt[0]), .Y(n1046) );
  NOR4X1 U784 ( .A(outpos[2]), .B(outpos[3]), .C(outpos[4]), .D(outpos[5]), 
        .Y(n1045) );
  XNOR2X1 U785 ( .A(n94), .B(n1048), .Y(\col_t[2] ) );
  OAI21XL U786 ( .A0(n385), .A1(n1049), .B0(n1050), .Y(n1048) );
  OAI2BB1X1 U787 ( .A0N(n1049), .A1N(n385), .B0(cnt[1]), .Y(n1050) );
  XNOR2X1 U788 ( .A(cnt[1]), .B(n385), .Y(n1051) );
  OR2X1 U789 ( .A(n386), .B(n96), .Y(n1049) );
  XNOR2X1 U790 ( .A(row[0]), .B(n93), .Y(N449) );
endmodule

