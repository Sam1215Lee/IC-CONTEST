
module JAM_DW01_add_0 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [9:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  AND2X2 U2 ( .A(A[7]), .B(carry[7]), .Y(n2) );
  XOR2XL U3 ( .A(A[8]), .B(n2), .Y(SUM[8]) );
  XNOR2X1 U4 ( .A(A[9]), .B(n3), .Y(SUM[9]) );
  XOR2XL U5 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U6 ( .A(A[8]), .B(n2), .Y(n3) );
  XOR2X1 U7 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
endmodule


module JAM_DW01_add_1 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3;
  wire   [9:1] carry;

  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  XOR2X1 U1 ( .A(n1), .B(A[9]), .Y(SUM[9]) );
  XOR2X1 U2 ( .A(A[8]), .B(n3), .Y(SUM[8]) );
  AND2X2 U3 ( .A(n3), .B(A[8]), .Y(n1) );
  AND2X2 U4 ( .A(B[0]), .B(A[0]), .Y(n2) );
  AND2XL U5 ( .A(A[7]), .B(carry[7]), .Y(n3) );
  XOR2XL U6 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2XL U7 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
endmodule


module JAM ( CLK, RST, W, J, Cost, MatchCount, MinCost, Valid );
  output [2:0] W;
  output [2:0] J;
  input [6:0] Cost;
  output [3:0] MatchCount;
  output [9:0] MinCost;
  input CLK, RST;
  output Valid;
  wire   N154, N155, N156, N157, N158, N159, N160, N161, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, \buff[7][2] , \buff[7][1] , \buff[7][0] , \buff[6][2] ,
         \buff[6][1] , \buff[6][0] , \buff[5][2] , \buff[5][1] , \buff[5][0] ,
         \buff[4][2] , \buff[4][1] , \buff[4][0] , \buff[3][2] , \buff[3][1] ,
         \buff[3][0] , \buff[2][2] , \buff[2][1] , \buff[2][0] , \buff[1][2] ,
         \buff[1][1] , \buff[1][0] , \buff[0][2] , \buff[0][1] , \buff[0][0] ,
         N180, N181, N183, N184, N185, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, \val[2] , N251, N252, N253, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N451, N452, n36, n38, n40,
         n41, n42, n46, n47, n49, n50, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n68, n69, n72, n73, n74, n76, n79, n81,
         n82, n83, n84, n86, n88, n89, n90, n91, n93, n95, n96, n97, n98, n99,
         n100, n102, n103, n105, n107, n108, n109, n110, n112, n113, n114,
         n116, n117, n121, n122, n123, n127, n129, n130, n131, n132, n133,
         n134, n135, n137, n139, n140, n141, n142, n143, n144, n145, n146,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n158, n159,
         n160, n161, n162, n163, n164, n165, n167, n168, n169, n170, n171,
         n172, n173, n175, n176, n177, n179, n180, n181, n182, n183, n184,
         n186, n187, n188, n189, n190, n191, n194, n195, n196, n198, n199,
         n200, n203, n204, n207, n209, n210, n211, n213, n214, n215, n217,
         n219, n220, n221, n222, n223, n225, n226, n227, n228, n230, n231,
         n232, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n246, n247, n248, n249, n250, n251, n252, n254, n255, n256, n258,
         n259, n262, n263, n264, n266, n267, n268, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n406, n408, n421,
         n423, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544;
  wire   [1:0] state;
  wire   [1:0] next;
  wire   [9:0] sum;

  JAM_DW01_add_0 add_159 ( .A(sum), .B({1'b0, 1'b0, 1'b0, Cost}), .CI(1'b0), 
        .SUM({N439, N438, N437, N436, N435, N434, N433, N432, N431, N430}) );
  JAM_DW01_add_1 add_86 ( .A({MinCost[9], n553, n554, n555, MinCost[5:3], n559, 
        n560, n561}), .B({1'b0, 1'b0, 1'b0, Cost}), .CI(1'b0), .SUM({N203, 
        N202, N201, N200, N199, N198, N197, N196, N195, N194}) );
  DFFQX1 \val_reg[2]  ( .D(n384), .CK(CLK), .Q(\val[2] ) );
  DFFX1 \val_reg[0]  ( .D(n386), .CK(CLK), .Q(n279), .QN(n541) );
  DFFSX1 \buff_reg[3][0]  ( .D(n369), .CK(CLK), .SN(n498), .Q(\buff[3][0] ), 
        .QN(n321) );
  DFFSX1 \buff_reg[7][0]  ( .D(n357), .CK(CLK), .SN(n446), .Q(\buff[7][0] ), 
        .QN(n291) );
  DFFX1 \val_reg[1]  ( .D(n385), .CK(CLK), .Q(n280), .QN(n540) );
  DFFRX1 cnt_reg ( .D(n391), .CK(CLK), .RN(n444), .QN(n309) );
  DFFRX1 \cur_reg[0]  ( .D(next[0]), .CK(CLK), .RN(n444), .Q(n400), .QN(n317)
         );
  DFFRX1 \buff_reg[3][2]  ( .D(n367), .CK(CLK), .RN(n445), .Q(\buff[3][2] ), 
        .QN(n284) );
  DFFRX1 \buff_reg[1][2]  ( .D(n373), .CK(CLK), .RN(n444), .Q(\buff[1][2] ), 
        .QN(n323) );
  DFFRX1 \buff_reg[1][1]  ( .D(n374), .CK(CLK), .RN(n444), .Q(\buff[1][1] ), 
        .QN(n324) );
  DFFRX1 \buff_reg[5][1]  ( .D(n362), .CK(CLK), .RN(n445), .Q(\buff[5][1] ), 
        .QN(n287) );
  DFFRX1 \buff_reg[0][2]  ( .D(n376), .CK(CLK), .RN(n444), .Q(\buff[0][2] ), 
        .QN(n326) );
  DFFRX1 \buff_reg[0][1]  ( .D(n377), .CK(CLK), .RN(n445), .Q(\buff[0][1] ), 
        .QN(n327) );
  DFFRX1 \buff_reg[0][0]  ( .D(n378), .CK(CLK), .RN(n444), .Q(\buff[0][0] ), 
        .QN(n328) );
  DFFRX1 \buff_reg[4][1]  ( .D(n365), .CK(CLK), .RN(n445), .Q(\buff[4][1] ), 
        .QN(n285) );
  DFFRX1 \buff_reg[4][0]  ( .D(n366), .CK(CLK), .RN(n445), .Q(\buff[4][0] ), 
        .QN(n320) );
  DFFRX1 \buff_reg[2][2]  ( .D(n370), .CK(CLK), .RN(n445), .Q(\buff[2][2] ), 
        .QN(n282) );
  DFFRX1 \buff_reg[2][0]  ( .D(n372), .CK(CLK), .RN(n445), .Q(\buff[2][0] ), 
        .QN(n322) );
  DFFRX1 \buff_reg[6][0]  ( .D(n360), .CK(CLK), .RN(n445), .Q(\buff[6][0] ), 
        .QN(n318) );
  DFFSX1 \buff_reg[3][1]  ( .D(n368), .CK(CLK), .SN(n498), .Q(\buff[3][1] ), 
        .QN(n283) );
  DFFSX1 \buff_reg[7][1]  ( .D(n356), .CK(CLK), .SN(n446), .Q(\buff[7][1] ), 
        .QN(n292) );
  DFFSX1 \buff_reg[7][2]  ( .D(n396), .CK(CLK), .SN(n446), .Q(\buff[7][2] ), 
        .QN(n293) );
  DFFSX1 \buff_reg[1][0]  ( .D(n375), .CK(CLK), .SN(n446), .Q(\buff[1][0] ), 
        .QN(n325) );
  DFFSX1 \buff_reg[5][0]  ( .D(n363), .CK(CLK), .SN(n446), .Q(\buff[5][0] ), 
        .QN(n319) );
  DFFSX1 \buff_reg[5][2]  ( .D(n361), .CK(CLK), .SN(n446), .Q(\buff[5][2] ), 
        .QN(n288) );
  DFFSX1 \buff_reg[4][2]  ( .D(n364), .CK(CLK), .SN(n446), .Q(\buff[4][2] ), 
        .QN(n286) );
  DFFSX1 \buff_reg[2][1]  ( .D(n371), .CK(CLK), .SN(n498), .Q(\buff[2][1] ), 
        .QN(n281) );
  DFFSX1 \buff_reg[6][2]  ( .D(n358), .CK(CLK), .SN(n498), .Q(\buff[6][2] ), 
        .QN(n290) );
  DFFSX1 \buff_reg[6][1]  ( .D(n359), .CK(CLK), .SN(n498), .Q(\buff[6][1] ), 
        .QN(n289) );
  DFFRX1 \state_reg[1]  ( .D(n388), .CK(CLK), .RN(n444), .Q(state[1]), .QN(
        n399) );
  DFFQX1 \sum_reg[5]  ( .D(n349), .CK(CLK), .Q(sum[5]) );
  DFFQX1 \sum_reg[6]  ( .D(n348), .CK(CLK), .Q(sum[6]) );
  DFFQX1 \sum_reg[4]  ( .D(n350), .CK(CLK), .Q(sum[4]) );
  DFFQX1 \sum_reg[3]  ( .D(n351), .CK(CLK), .Q(sum[3]) );
  DFFQX1 \sum_reg[2]  ( .D(n352), .CK(CLK), .Q(sum[2]) );
  DFFRX1 \sub1_reg[1]  ( .D(n381), .CK(CLK), .RN(n444), .Q(N157), .QN(n334) );
  DFFQX1 \sum_reg[7]  ( .D(n347), .CK(CLK), .Q(sum[7]) );
  DFFQX1 \sum_reg[1]  ( .D(n353), .CK(CLK), .Q(sum[1]) );
  DFFQX1 \sum_reg[0]  ( .D(n354), .CK(CLK), .Q(sum[0]) );
  DFFRX1 \cur_reg[1]  ( .D(next[1]), .CK(CLK), .RN(n444), .QN(n316) );
  DFFQX1 \sum_reg[9]  ( .D(n355), .CK(CLK), .Q(sum[9]) );
  DFFQX1 \sum_reg[8]  ( .D(n346), .CK(CLK), .Q(sum[8]) );
  DFFRX1 \MinCost_reg[3]  ( .D(n493), .CK(CLK), .RN(n446), .Q(n558), .QN(n423)
         );
  DFFRX1 \MinCost_reg[4]  ( .D(n492), .CK(CLK), .RN(n446), .Q(n557), .QN(n421)
         );
  DFFRX1 \MinCost_reg[0]  ( .D(n496), .CK(CLK), .RN(n445), .Q(n561), .QN(n426)
         );
  DFFRX1 \MinCost_reg[6]  ( .D(n490), .CK(CLK), .RN(n445), .Q(n555), .QN(n479)
         );
  DFFRX1 \MinCost_reg[2]  ( .D(n494), .CK(CLK), .RN(n446), .Q(n559), .QN(n430)
         );
  DFFQX1 Valid_reg ( .D(n297), .CK(CLK), .Q(n562) );
  DFFSX1 \W_reg[0]  ( .D(n393), .CK(CLK), .SN(n446), .Q(n548), .QN(n315) );
  DFFSX1 \W_reg[1]  ( .D(n392), .CK(CLK), .SN(n446), .Q(n547), .QN(n314) );
  DFFSX1 \J_reg[0]  ( .D(n345), .CK(CLK), .SN(n446), .Q(n550), .QN(n332) );
  DFFSX1 \J_reg[2]  ( .D(n343), .CK(CLK), .SN(n446), .Q(n549), .QN(n294) );
  DFFRX1 \MatchCount_reg[3]  ( .D(n339), .CK(CLK), .RN(n446), .Q(n551), .QN(
        n329) );
  DFFRX1 \MatchCount_reg[1]  ( .D(n341), .CK(CLK), .RN(n446), .Q(n552), .QN(
        n296) );
  DFFRX1 \MatchCount_reg[2]  ( .D(n340), .CK(CLK), .RN(n446), .QN(n330) );
  DFFRX1 \MinCost_reg[1]  ( .D(n495), .CK(CLK), .RN(n446), .Q(n560), .QN(n408)
         );
  DFFRX1 \MinCost_reg[5]  ( .D(n491), .CK(CLK), .RN(n445), .Q(n556), .QN(n406)
         );
  DFFRX1 \MatchCount_reg[0]  ( .D(n342), .CK(CLK), .RN(n446), .QN(n295) );
  DFFRX1 \sub1_reg[2]  ( .D(n383), .CK(CLK), .RN(n498), .Q(N158), .QN(n333) );
  DFFRX1 \MinCost_reg[7]  ( .D(n489), .CK(CLK), .RN(n498), .Q(n554), .QN(n480)
         );
  DFFSXL \J_reg[1]  ( .D(n344), .CK(CLK), .SN(n498), .Q(n544), .QN(n331) );
  DFFRX2 \sub1_reg[0]  ( .D(n382), .CK(CLK), .RN(n498), .Q(N156), .QN(n335) );
  DFFRX1 \state_reg[0]  ( .D(n387), .CK(CLK), .RN(n498), .Q(state[0]), .QN(
        n530) );
  DFFSX4 \index_reg[0]  ( .D(n390), .CK(CLK), .SN(n498), .Q(n531), .QN(n312)
         );
  DFFSX2 \index_reg[2]  ( .D(n395), .CK(CLK), .SN(n498), .Q(N155), .QN(n310)
         );
  DFFSX4 \index_reg[1]  ( .D(n389), .CK(CLK), .SN(n498), .Q(N154), .QN(n311)
         );
  DFFSX2 \sub2_reg[0]  ( .D(n397), .CK(CLK), .SN(n498), .Q(N159), .QN(n338) );
  DFFSX2 \sub2_reg[1]  ( .D(n380), .CK(CLK), .SN(n498), .Q(N160), .QN(n337) );
  DFFSX2 \sub2_reg[2]  ( .D(n379), .CK(CLK), .SN(n498), .Q(N161), .QN(n336) );
  DFFSX1 \W_reg[2]  ( .D(n394), .CK(CLK), .SN(n498), .QN(n313) );
  DFFRX1 \MinCost_reg[8]  ( .D(n488), .CK(CLK), .RN(n445), .Q(n553) );
  DFFRX1 \MinCost_reg[9]  ( .D(n487), .CK(CLK), .RN(n445), .QN(n401) );
  AOI222X1 U322 ( .A0(N203), .A1(n538), .B0(sum[9]), .B1(n52), .C0(n443), .C1(
        MinCost[9]), .Y(n54) );
  CLKINVX1 U323 ( .A(n62), .Y(n488) );
  AOI222X1 U324 ( .A0(N202), .A1(n538), .B0(sum[8]), .B1(n52), .C0(n443), .C1(
        MinCost[8]), .Y(n62) );
  CLKINVX1 U325 ( .A(n54), .Y(n487) );
  INVX16 U326 ( .A(n401), .Y(MinCost[9]) );
  CLKMX2X2 U327 ( .A(n447), .B(n448), .S0(N155), .Y(n398) );
  CLKBUFX2 U328 ( .A(n445), .Y(n444) );
  INVX3 U329 ( .A(RST), .Y(n498) );
  CLKINVX1 U330 ( .A(n544), .Y(n402) );
  INVX16 U331 ( .A(n402), .Y(J[1]) );
  INVX16 U332 ( .A(n313), .Y(W[2]) );
  OAI22X1 U333 ( .A0(sum[9]), .A1(n401), .B0(n486), .B1(n472), .Y(N451) );
  INVX16 U334 ( .A(n295), .Y(MatchCount[0]) );
  INVX16 U335 ( .A(n406), .Y(MinCost[5]) );
  INVX12 U336 ( .A(n408), .Y(MinCost[1]) );
  AO21XL U337 ( .A0(n485), .A1(n462), .B0(n560), .Y(n461) );
  INVX16 U338 ( .A(n330), .Y(MatchCount[2]) );
  BUFX12 U339 ( .A(n552), .Y(MatchCount[1]) );
  BUFX12 U340 ( .A(n551), .Y(MatchCount[3]) );
  BUFX12 U341 ( .A(n549), .Y(J[2]) );
  BUFX12 U342 ( .A(n550), .Y(J[0]) );
  BUFX12 U343 ( .A(n547), .Y(W[1]) );
  BUFX12 U344 ( .A(n548), .Y(W[0]) );
  BUFX16 U345 ( .A(n562), .Y(Valid) );
  BUFX12 U346 ( .A(n559), .Y(MinCost[2]) );
  INVX12 U347 ( .A(n479), .Y(MinCost[6]) );
  BUFX12 U348 ( .A(n561), .Y(MinCost[0]) );
  INVX12 U349 ( .A(n480), .Y(MinCost[7]) );
  INVX16 U350 ( .A(n421), .Y(MinCost[4]) );
  NOR2XL U351 ( .A(n484), .B(n557), .Y(n475) );
  INVX16 U352 ( .A(n423), .Y(MinCost[3]) );
  NOR2BXL U353 ( .AN(sum[3]), .B(n558), .Y(n476) );
  BUFX12 U354 ( .A(n553), .Y(MinCost[8]) );
  AOI32XL U355 ( .A0(n471), .A1(n482), .A2(n470), .B0(n553), .B1(n481), .Y(
        n472) );
  INVX1 U356 ( .A(n74), .Y(n533) );
  NOR2X1 U357 ( .A(n426), .B(sum[0]), .Y(n462) );
  AOI2BB1X1 U358 ( .A0N(n41), .A1N(n543), .B0(n538), .Y(n53) );
  OAI222XL U359 ( .A0(n469), .A1(n468), .B0(sum[6]), .B1(n479), .C0(sum[7]), 
        .C1(n480), .Y(n470) );
  NAND2BX1 U360 ( .AN(n467), .B(n466), .Y(n468) );
  BUFX2 U361 ( .A(n53), .Y(n443) );
  NOR2XL U362 ( .A(n483), .B(n556), .Y(n467) );
  OAI21XL U363 ( .A0(n329), .A1(n63), .B0(n64), .Y(n339) );
  NOR2XL U364 ( .A(n481), .B(n553), .Y(n460) );
  AND2XL U365 ( .A(n556), .B(n483), .Y(n427) );
  AND2XL U366 ( .A(n557), .B(n484), .Y(n428) );
  AND2X2 U367 ( .A(n465), .B(n464), .Y(n429) );
  NOR3X1 U368 ( .A(n427), .B(n428), .C(n429), .Y(n469) );
  NOR2X1 U369 ( .A(n476), .B(n475), .Y(n465) );
  OR2X1 U370 ( .A(n534), .B(n68), .Y(n431) );
  NAND2X1 U371 ( .A(n431), .B(n443), .Y(n74) );
  NAND2X1 U372 ( .A(n432), .B(n532), .Y(n69) );
  NAND3BXL U373 ( .AN(N451), .B(n474), .C(n473), .Y(n477) );
  OAI21X1 U374 ( .A0(n268), .A1(n529), .B0(n528), .Y(n183) );
  OAI21X1 U375 ( .A0(n210), .A1(n211), .B0(n38), .Y(n184) );
  NOR2X1 U376 ( .A(n399), .B(n530), .Y(n267) );
  NAND3X1 U377 ( .A(n535), .B(n38), .C(n83), .Y(n89) );
  INVX1 U378 ( .A(n65), .Y(n532) );
  OA21XL U379 ( .A0(MatchCount[2]), .A1(n68), .B0(n69), .Y(n63) );
  OA21XL U380 ( .A0(MatchCount[0]), .A1(n68), .B0(n74), .Y(n72) );
  NOR2BXL U381 ( .AN(sum[0]), .B(n561), .Y(n457) );
  AOI32X1 U382 ( .A0(n270), .A1(n196), .A2(n271), .B0(N155), .B1(n333), .Y(
        n268) );
  NOR4X1 U383 ( .A(n315), .B(n314), .C(n313), .D(n309), .Y(n36) );
  NOR2X1 U384 ( .A(n399), .B(state[0]), .Y(n181) );
  NAND2X1 U385 ( .A(n316), .B(n400), .Y(n91) );
  OA21XL U386 ( .A0(n334), .A1(N156), .B0(n135), .Y(n187) );
  NOR2X1 U387 ( .A(state[0]), .B(state[1]), .Y(n198) );
  NAND3X1 U388 ( .A(state[0]), .B(n399), .C(n537), .Y(n211) );
  NAND3X1 U389 ( .A(N160), .B(N161), .C(n338), .Y(n112) );
  NAND3X1 U390 ( .A(n338), .B(N160), .C(n336), .Y(n161) );
  NAND3X1 U391 ( .A(n338), .B(N161), .C(n337), .Y(n142) );
  NAND3X1 U392 ( .A(N159), .B(N161), .C(n337), .Y(n132) );
  NAND3X1 U393 ( .A(N159), .B(N160), .C(n336), .Y(n151) );
  NAND3X1 U394 ( .A(n337), .B(N159), .C(n336), .Y(n170) );
  NAND3X1 U395 ( .A(n337), .B(n338), .C(n336), .Y(n176) );
  NAND4XL U396 ( .A(n296), .B(n536), .C(n74), .D(MatchCount[0]), .Y(n73) );
  OR2XL U397 ( .A(n536), .B(n533), .Y(n432) );
  INVXL U398 ( .A(n68), .Y(n536) );
  NOR2X2 U399 ( .A(n535), .B(n443), .Y(n52) );
  CLKINVX1 U400 ( .A(n203), .Y(n497) );
  OAI221XL U401 ( .A0(n509), .A1(n47), .B0(n522), .B1(n535), .C0(n239), .Y(
        n227) );
  NOR2BX1 U402 ( .AN(n41), .B(n240), .Y(n239) );
  NAND3X2 U403 ( .A(n267), .B(n517), .C(n537), .Y(n121) );
  CLKINVX1 U404 ( .A(n137), .Y(n503) );
  CLKINVX1 U405 ( .A(n127), .Y(n499) );
  CLKINVX1 U406 ( .A(n146), .Y(n500) );
  CLKINVX1 U407 ( .A(n165), .Y(n501) );
  NAND2BX1 U408 ( .AN(n199), .B(n200), .Y(n191) );
  NAND2X1 U409 ( .A(n102), .B(n266), .Y(n99) );
  CLKINVX1 U410 ( .A(n221), .Y(n514) );
  OAI2BB1X1 U411 ( .A0N(n266), .A1N(n529), .B0(n102), .Y(n100) );
  CLKINVX1 U412 ( .A(n173), .Y(n505) );
  NOR2BX1 U413 ( .AN(n38), .B(n227), .Y(n223) );
  NAND2X1 U414 ( .A(n191), .B(n183), .Y(n188) );
  NOR3X1 U415 ( .A(n509), .B(n209), .C(n47), .Y(n199) );
  NAND2X1 U416 ( .A(n267), .B(n184), .Y(n186) );
  CLKINVX1 U417 ( .A(n184), .Y(n510) );
  CLKINVX1 U418 ( .A(n215), .Y(n509) );
  INVX3 U419 ( .A(n267), .Y(n529) );
  CLKINVX1 U420 ( .A(n89), .Y(n518) );
  NOR2X2 U421 ( .A(n524), .B(n529), .Y(n114) );
  NOR2X2 U422 ( .A(n523), .B(n529), .Y(n108) );
  NAND2X1 U423 ( .A(n537), .B(n89), .Y(n231) );
  INVX3 U424 ( .A(n240), .Y(n527) );
  CLKINVX1 U425 ( .A(n214), .Y(n516) );
  OA21XL U426 ( .A0(n209), .A1(n47), .B0(n200), .Y(n220) );
  CLKINVX1 U427 ( .A(n209), .Y(n522) );
  INVXL U428 ( .A(N451), .Y(n543) );
  NAND3X1 U429 ( .A(n79), .B(n543), .C(N452), .Y(n68) );
  OAI21X1 U430 ( .A0(n207), .A1(n199), .B0(n444), .Y(n203) );
  NOR2X1 U431 ( .A(n210), .B(n211), .Y(n207) );
  OAI221XL U432 ( .A0(n497), .A1(n539), .B0(n523), .B1(n203), .C0(n204), .Y(
        n384) );
  NAND2X1 U433 ( .A(n497), .B(n198), .Y(n204) );
  CLKBUFX3 U434 ( .A(n96), .Y(n442) );
  NOR2X1 U435 ( .A(n95), .B(n535), .Y(n96) );
  OAI222X4 U436 ( .A0(n266), .A1(n527), .B0(n123), .B1(n154), .C0(n121), .C1(
        n250), .Y(n102) );
  OAI222X1 U437 ( .A0(n121), .A1(n140), .B0(n527), .B1(n142), .C0(n123), .C1(
        n145), .Y(n137) );
  OAI222X1 U438 ( .A0(n121), .A1(n130), .B0(n527), .B1(n132), .C0(n123), .C1(
        n135), .Y(n127) );
  OAI222X1 U439 ( .A0(n527), .A1(n151), .B0(n154), .B1(n155), .C0(n121), .C1(
        n149), .Y(n146) );
  OAI222X1 U440 ( .A0(n135), .A1(n155), .B0(n527), .B1(n170), .C0(n121), .C1(
        n168), .Y(n165) );
  OAI211X1 U441 ( .A0(n515), .A1(n211), .B0(n535), .C0(n220), .Y(n221) );
  CLKINVX1 U442 ( .A(n219), .Y(n515) );
  OAI22X1 U443 ( .A0(n527), .A1(n176), .B0(n145), .B1(n155), .Y(n173) );
  OAI211X1 U444 ( .A0(n523), .A1(n241), .B0(n242), .C0(n243), .Y(n215) );
  OAI211X1 U445 ( .A0(N180), .A1(n512), .B0(N181), .C0(n513), .Y(n243) );
  OAI221XL U446 ( .A0(N181), .A1(n513), .B0(N180), .B1(n512), .C0(n246), .Y(
        n242) );
  CLKINVX1 U447 ( .A(n251), .Y(n513) );
  NAND3X1 U448 ( .A(n267), .B(n268), .C(n537), .Y(n38) );
  INVX3 U449 ( .A(N181), .Y(n524) );
  CLKINVX1 U450 ( .A(n105), .Y(n502) );
  CLKINVX1 U451 ( .A(n156), .Y(n504) );
  CLKINVX1 U452 ( .A(N180), .Y(n523) );
  NAND2X1 U453 ( .A(N156), .B(n542), .Y(n154) );
  CLKINVX1 U454 ( .A(n268), .Y(n517) );
  OAI22XL U455 ( .A0(N180), .A1(n525), .B0(n277), .B1(n278), .Y(n276) );
  NOR2X1 U456 ( .A(n441), .B(n524), .Y(n278) );
  AOI211X1 U457 ( .A0(n441), .A1(n524), .B0(n398), .C0(N185), .Y(n277) );
  NAND3X1 U458 ( .A(N154), .B(N155), .C(n531), .Y(n250) );
  NAND2X1 U459 ( .A(n198), .B(n191), .Y(n190) );
  OAI2BB1X1 U460 ( .A0N(N155), .A1N(n194), .B0(n262), .Y(n219) );
  AOI33X1 U461 ( .A0(n263), .A1(N154), .A2(n187), .B0(N156), .B1(n531), .B2(
        n264), .Y(n262) );
  OA21XL U462 ( .A0(n187), .A1(N154), .B0(n263), .Y(n264) );
  OR2X1 U463 ( .A(n194), .B(N155), .Y(n263) );
  INVX3 U464 ( .A(n181), .Y(n528) );
  CLKINVX1 U465 ( .A(n241), .Y(n512) );
  CLKINVX1 U466 ( .A(N183), .Y(n525) );
  NOR2X2 U467 ( .A(n398), .B(n529), .Y(n117) );
  OAI22X1 U468 ( .A0(n529), .A1(n140), .B0(n528), .B1(n142), .Y(n141) );
  OAI22X1 U469 ( .A0(n529), .A1(n159), .B0(n528), .B1(n161), .Y(n160) );
  OAI22X1 U470 ( .A0(n529), .A1(n168), .B0(n528), .B1(n170), .Y(n169) );
  OAI22X1 U471 ( .A0(n529), .A1(n149), .B0(n528), .B1(n151), .Y(n150) );
  OAI22X1 U472 ( .A0(n529), .A1(n109), .B0(n528), .B1(n112), .Y(n110) );
  OAI22X1 U473 ( .A0(n529), .A1(n130), .B0(n528), .B1(n132), .Y(n131) );
  NAND2X1 U474 ( .A(n198), .B(n537), .Y(n47) );
  OAI21X1 U475 ( .A0(n211), .A1(n219), .B0(n220), .Y(n214) );
  CLKINVX1 U476 ( .A(n98), .Y(n507) );
  CLKINVX1 U477 ( .A(n179), .Y(n506) );
  CLKINVX1 U478 ( .A(n103), .Y(n508) );
  NOR2X1 U479 ( .A(n159), .B(N154), .Y(n209) );
  OAI211X1 U480 ( .A0(n36), .A1(n535), .B0(n38), .C0(n521), .Y(next[1]) );
  NAND2X1 U481 ( .A(n36), .B(n79), .Y(n41) );
  NOR2X1 U482 ( .A(n528), .B(n91), .Y(n240) );
  INVX3 U483 ( .A(n83), .Y(n538) );
  INVX3 U484 ( .A(n79), .Y(n535) );
  INVX3 U485 ( .A(n91), .Y(n537) );
  NAND3X1 U486 ( .A(N160), .B(N161), .C(N159), .Y(n266) );
  CLKINVX1 U487 ( .A(n36), .Y(n534) );
  NAND4X1 U488 ( .A(n521), .B(n40), .C(n41), .D(n42), .Y(next[0]) );
  OAI21XL U489 ( .A0(n517), .A1(n529), .B0(n537), .Y(n40) );
  OA21XL U490 ( .A0(n529), .A1(n91), .B0(n527), .Y(n200) );
  NOR2X1 U491 ( .A(n176), .B(n528), .Y(n177) );
  NOR2X1 U492 ( .A(J[1]), .B(n88), .Y(n86) );
  CLKBUFX3 U493 ( .A(n498), .Y(n446) );
  CLKBUFX3 U494 ( .A(n498), .Y(n445) );
  CLKINVX1 U495 ( .A(n474), .Y(n486) );
  CLKINVX1 U496 ( .A(n460), .Y(n482) );
  OAI32X1 U497 ( .A0(MatchCount[2]), .A1(n68), .A2(n532), .B0(n330), .B1(n69), 
        .Y(n340) );
  OAI22XL U498 ( .A0(n295), .A1(n74), .B0(n533), .B1(n76), .Y(n342) );
  NOR3XL U499 ( .A(n295), .B(N451), .C(n538), .Y(n76) );
  NOR3X1 U500 ( .A(n296), .B(n295), .C(n533), .Y(n65) );
  OAI21XL U501 ( .A0(n296), .A1(n72), .B0(n73), .Y(n341) );
  NAND4X1 U502 ( .A(n329), .B(n65), .C(n536), .D(MatchCount[2]), .Y(n64) );
  CLKINVX1 U503 ( .A(n50), .Y(n496) );
  AOI222XL U504 ( .A0(N194), .A1(n538), .B0(sum[0]), .B1(n52), .C0(n443), .C1(
        MinCost[0]), .Y(n50) );
  CLKINVX1 U505 ( .A(n61), .Y(n489) );
  AOI222XL U506 ( .A0(N201), .A1(n538), .B0(sum[7]), .B1(n52), .C0(n443), .C1(
        n554), .Y(n61) );
  CLKINVX1 U507 ( .A(n57), .Y(n493) );
  AOI222XL U508 ( .A0(N197), .A1(n538), .B0(sum[3]), .B1(n52), .C0(n443), .C1(
        MinCost[3]), .Y(n57) );
  CLKINVX1 U509 ( .A(n55), .Y(n495) );
  AOI222XL U510 ( .A0(N195), .A1(n538), .B0(sum[1]), .B1(n52), .C0(n443), .C1(
        MinCost[1]), .Y(n55) );
  CLKINVX1 U511 ( .A(n58), .Y(n492) );
  AOI222XL U512 ( .A0(N198), .A1(n538), .B0(sum[4]), .B1(n52), .C0(n443), .C1(
        MinCost[4]), .Y(n58) );
  CLKINVX1 U513 ( .A(n59), .Y(n491) );
  AOI222XL U514 ( .A0(N199), .A1(n538), .B0(sum[5]), .B1(n52), .C0(n443), .C1(
        MinCost[5]), .Y(n59) );
  CLKINVX1 U515 ( .A(n56), .Y(n494) );
  AOI222XL U516 ( .A0(N196), .A1(n538), .B0(sum[2]), .B1(n52), .C0(n443), .C1(
        MinCost[2]), .Y(n56) );
  CLKINVX1 U517 ( .A(n60), .Y(n490) );
  AOI222XL U518 ( .A0(N200), .A1(n538), .B0(sum[6]), .B1(n52), .C0(n443), .C1(
        n555), .Y(n60) );
  AO22X1 U519 ( .A0(n95), .A1(sum[9]), .B0(N439), .B1(n442), .Y(n355) );
  AO22X1 U520 ( .A0(n95), .A1(sum[8]), .B0(N438), .B1(n442), .Y(n346) );
  AO22X1 U521 ( .A0(n95), .A1(sum[7]), .B0(N437), .B1(n442), .Y(n347) );
  OAI221XL U522 ( .A0(n497), .A1(n540), .B0(n524), .B1(n203), .C0(n204), .Y(
        n385) );
  OAI221XL U523 ( .A0(n497), .A1(n541), .B0(n398), .B1(n203), .C0(n204), .Y(
        n386) );
  NAND2X2 U524 ( .A(n444), .B(n97), .Y(n95) );
  OAI2BB1X1 U525 ( .A0N(n79), .A1N(n309), .B0(n38), .Y(n97) );
  CLKINVX1 U526 ( .A(sum[1]), .Y(n485) );
  CLKINVX1 U527 ( .A(sum[4]), .Y(n484) );
  AO22X1 U528 ( .A0(n95), .A1(sum[0]), .B0(N430), .B1(n442), .Y(n354) );
  AO22X1 U529 ( .A0(n95), .A1(sum[6]), .B0(N436), .B1(n442), .Y(n348) );
  AO22X1 U530 ( .A0(n95), .A1(sum[5]), .B0(N435), .B1(n442), .Y(n349) );
  AO22X1 U531 ( .A0(n95), .A1(sum[4]), .B0(N434), .B1(n442), .Y(n350) );
  AO22X1 U532 ( .A0(n95), .A1(sum[3]), .B0(N433), .B1(n442), .Y(n351) );
  AO22X1 U533 ( .A0(n95), .A1(sum[2]), .B0(N432), .B1(n442), .Y(n352) );
  AO22X1 U534 ( .A0(n95), .A1(sum[1]), .B0(N431), .B1(n442), .Y(n353) );
  XOR2XL U535 ( .A(Valid), .B(n49), .Y(n297) );
  NOR3X1 U536 ( .A(RST), .B(n316), .C(n317), .Y(n49) );
  CLKINVX1 U537 ( .A(sum[5]), .Y(n483) );
  CLKINVX1 U538 ( .A(sum[8]), .Y(n481) );
  OAI221X1 U539 ( .A0(n527), .A1(n112), .B0(n121), .B1(n109), .C0(n122), .Y(
        n105) );
  NAND3BX1 U540 ( .AN(n123), .B(n335), .C(n542), .Y(n122) );
  OAI221X1 U541 ( .A0(n527), .A1(n161), .B0(n159), .B1(n121), .C0(n164), .Y(
        n156) );
  NAND3BX1 U542 ( .AN(n155), .B(n335), .C(n542), .Y(n164) );
  AOI2BB2X1 U543 ( .B0(n542), .B1(n312), .A0N(n333), .A1N(N155), .Y(n270) );
  OAI2BB1X1 U544 ( .A0N(n154), .A1N(N154), .B0(n145), .Y(n271) );
  CLKMX2X2 U545 ( .A(n433), .B(n434), .S0(N155), .Y(N180) );
  MX4X1 U546 ( .A(\buff[0][2] ), .B(\buff[1][2] ), .C(\buff[2][2] ), .D(
        \buff[3][2] ), .S0(n531), .S1(N154), .Y(n433) );
  MX4X1 U547 ( .A(\buff[4][2] ), .B(\buff[5][2] ), .C(\buff[6][2] ), .D(
        \buff[7][2] ), .S0(n531), .S1(N154), .Y(n434) );
  OAI211X1 U548 ( .A0(\val[2] ), .A1(n523), .B0(n272), .C0(n273), .Y(n210) );
  OAI22XL U549 ( .A0(n274), .A1(n275), .B0(N180), .B1(n539), .Y(n273) );
  OAI21XL U550 ( .A0(N183), .A1(n523), .B0(n276), .Y(n272) );
  NOR2X1 U551 ( .A(n280), .B(n524), .Y(n275) );
  NAND2X2 U552 ( .A(n310), .B(n311), .Y(n168) );
  OAI222XL U553 ( .A0(n99), .A1(n103), .B0(n100), .B1(n511), .C0(n291), .C1(
        n102), .Y(n357) );
  CLKINVX1 U554 ( .A(N185), .Y(n511) );
  OAI222XL U555 ( .A0(n98), .A1(n99), .B0(n100), .B1(n526), .C0(n292), .C1(
        n102), .Y(n356) );
  CLKINVX1 U556 ( .A(n441), .Y(n526) );
  OAI222XL U557 ( .A0(n99), .A1(n179), .B0(n100), .B1(n525), .C0(n293), .C1(
        n102), .Y(n396) );
  OAI222XL U558 ( .A0(n187), .A1(n188), .B0(n189), .B1(n190), .C0(n334), .C1(
        n191), .Y(n381) );
  OAI222XL U559 ( .A0(n188), .A1(n194), .B0(n190), .B1(n195), .C0(n333), .C1(
        n191), .Y(n383) );
  NAND2X1 U560 ( .A(n196), .B(N155), .Y(n195) );
  OAI222XL U561 ( .A0(N156), .A1(n188), .B0(n531), .B1(n190), .C0(n335), .C1(
        n191), .Y(n382) );
  NAND3X2 U562 ( .A(n531), .B(N154), .C(n310), .Y(n149) );
  NAND3X2 U563 ( .A(N154), .B(N155), .C(n312), .Y(n109) );
  NAND3X2 U564 ( .A(n531), .B(N155), .C(n311), .Y(n130) );
  CLKMX2X2 U565 ( .A(n435), .B(n436), .S0(N155), .Y(N181) );
  MX4X1 U566 ( .A(\buff[0][1] ), .B(\buff[1][1] ), .C(\buff[2][1] ), .D(
        \buff[3][1] ), .S0(n531), .S1(N154), .Y(n435) );
  MX4X1 U567 ( .A(\buff[4][1] ), .B(\buff[5][1] ), .C(\buff[6][1] ), .D(
        \buff[7][1] ), .S0(n531), .S1(N154), .Y(n436) );
  CLKMX2X2 U568 ( .A(n437), .B(n438), .S0(N158), .Y(N183) );
  MX4X1 U569 ( .A(\buff[0][2] ), .B(\buff[1][2] ), .C(\buff[2][2] ), .D(
        \buff[3][2] ), .S0(N156), .S1(N157), .Y(n437) );
  MX4X1 U570 ( .A(\buff[4][2] ), .B(\buff[5][2] ), .C(\buff[6][2] ), .D(
        \buff[7][2] ), .S0(N156), .S1(N157), .Y(n438) );
  AOI211X1 U571 ( .A0(n280), .A1(n524), .B0(n398), .C0(n279), .Y(n274) );
  XNOR2X1 U572 ( .A(n333), .B(n154), .Y(n194) );
  CLKMX2X2 U573 ( .A(n439), .B(n440), .S0(N158), .Y(N185) );
  MX4X1 U574 ( .A(\buff[0][0] ), .B(\buff[1][0] ), .C(\buff[2][0] ), .D(
        \buff[3][0] ), .S0(N156), .S1(N157), .Y(n439) );
  MX4X1 U575 ( .A(\buff[4][0] ), .B(\buff[5][0] ), .C(\buff[6][0] ), .D(
        \buff[7][0] ), .S0(N156), .S1(N157), .Y(n440) );
  OAI221XL U576 ( .A0(n338), .A1(n184), .B0(n312), .B1(n510), .C0(n186), .Y(
        n397) );
  NAND2X1 U577 ( .A(n311), .B(n312), .Y(n196) );
  OAI221XL U578 ( .A0(n336), .A1(n184), .B0(n310), .B1(n510), .C0(n186), .Y(
        n379) );
  OAI221XL U579 ( .A0(n337), .A1(n184), .B0(n311), .B1(n510), .C0(n186), .Y(
        n380) );
  NAND2X2 U580 ( .A(n310), .B(n312), .Y(n159) );
  OAI31XL U581 ( .A0(n247), .A1(n248), .A2(n249), .B0(n398), .Y(n246) );
  OAI22XL U582 ( .A0(n325), .A1(n159), .B0(n328), .B1(n168), .Y(n248) );
  OAI22XL U583 ( .A0(n322), .A1(n149), .B0(n321), .B1(n140), .Y(n249) );
  OAI222XL U584 ( .A0(n320), .A1(n130), .B0(n319), .B1(n109), .C0(n318), .C1(
        n250), .Y(n247) );
  OAI211X1 U585 ( .A0(n83), .A1(n230), .B0(n231), .C0(n232), .Y(n392) );
  AOI2BB2X1 U586 ( .B0(n79), .B1(N154), .A0N(n234), .A1N(n314), .Y(n232) );
  OR2X2 U587 ( .A(n196), .B(n310), .Y(n140) );
  NAND3X1 U588 ( .A(n183), .B(N158), .C(n537), .Y(n123) );
  NAND3X1 U589 ( .A(n333), .B(n183), .C(n537), .Y(n155) );
  MXI4X1 U590 ( .A(\buff[0][0] ), .B(\buff[1][0] ), .C(\buff[2][0] ), .D(
        \buff[3][0] ), .S0(n531), .S1(N154), .Y(n447) );
  MXI4X1 U591 ( .A(\buff[4][0] ), .B(\buff[5][0] ), .C(\buff[6][0] ), .D(
        \buff[7][0] ), .S0(n531), .S1(N154), .Y(n448) );
  OAI22XL U592 ( .A0(n325), .A1(n165), .B0(n501), .B1(n172), .Y(n375) );
  AOI222XL U593 ( .A0(n117), .A1(n168), .B0(N185), .B1(n169), .C0(n508), .C1(
        n170), .Y(n172) );
  OAI22XL U594 ( .A0(n286), .A1(n137), .B0(n503), .B1(n139), .Y(n364) );
  AOI222XL U595 ( .A0(n108), .A1(n140), .B0(N183), .B1(n141), .C0(n506), .C1(
        n142), .Y(n139) );
  OAI22XL U596 ( .A0(n288), .A1(n127), .B0(n499), .B1(n129), .Y(n361) );
  AOI222XL U597 ( .A0(n108), .A1(n130), .B0(N183), .B1(n131), .C0(n506), .C1(
        n132), .Y(n129) );
  OAI22XL U598 ( .A0(n283), .A1(n146), .B0(n500), .B1(n152), .Y(n368) );
  AOI222XL U599 ( .A0(n114), .A1(n149), .B0(n441), .B1(n150), .C0(n507), .C1(
        n151), .Y(n152) );
  OAI22XL U600 ( .A0(n319), .A1(n127), .B0(n499), .B1(n134), .Y(n363) );
  AOI222XL U601 ( .A0(n117), .A1(n130), .B0(N185), .B1(n131), .C0(n508), .C1(
        n132), .Y(n134) );
  OAI22XL U602 ( .A0(n321), .A1(n146), .B0(n500), .B1(n153), .Y(n369) );
  AOI222XL U603 ( .A0(n117), .A1(n149), .B0(N185), .B1(n150), .C0(n508), .C1(
        n151), .Y(n153) );
  OAI22XL U604 ( .A0(n320), .A1(n137), .B0(n503), .B1(n144), .Y(n366) );
  AOI222XL U605 ( .A0(n117), .A1(n140), .B0(N185), .B1(n141), .C0(n508), .C1(
        n142), .Y(n144) );
  OAI22XL U606 ( .A0(n285), .A1(n137), .B0(n503), .B1(n143), .Y(n365) );
  AOI222XL U607 ( .A0(n114), .A1(n140), .B0(n441), .B1(n141), .C0(n507), .C1(
        n142), .Y(n143) );
  OAI22XL U608 ( .A0(n287), .A1(n127), .B0(n499), .B1(n133), .Y(n362) );
  AOI222XL U609 ( .A0(n114), .A1(n130), .B0(n441), .B1(n131), .C0(n507), .C1(
        n132), .Y(n133) );
  OAI22XL U610 ( .A0(n284), .A1(n146), .B0(n500), .B1(n148), .Y(n367) );
  AOI222XL U611 ( .A0(n108), .A1(n149), .B0(N183), .B1(n150), .C0(n506), .C1(
        n151), .Y(n148) );
  OAI22XL U612 ( .A0(n324), .A1(n165), .B0(n501), .B1(n171), .Y(n374) );
  AOI222XL U613 ( .A0(n114), .A1(n168), .B0(n441), .B1(n169), .C0(n507), .C1(
        n170), .Y(n171) );
  OAI22XL U614 ( .A0(n323), .A1(n165), .B0(n501), .B1(n167), .Y(n373) );
  AOI222XL U615 ( .A0(n108), .A1(n168), .B0(N183), .B1(n169), .C0(n506), .C1(
        n170), .Y(n167) );
  OAI22XL U616 ( .A0(n289), .A1(n105), .B0(n502), .B1(n113), .Y(n359) );
  AOI222XL U617 ( .A0(n114), .A1(n109), .B0(n441), .B1(n110), .C0(n507), .C1(
        n112), .Y(n113) );
  OAI22XL U618 ( .A0(n290), .A1(n105), .B0(n502), .B1(n107), .Y(n358) );
  AOI222XL U619 ( .A0(n108), .A1(n109), .B0(N183), .B1(n110), .C0(n506), .C1(
        n112), .Y(n107) );
  OAI22XL U620 ( .A0(n281), .A1(n156), .B0(n504), .B1(n162), .Y(n371) );
  AOI222XL U621 ( .A0(n114), .A1(n159), .B0(n441), .B1(n160), .C0(n507), .C1(
        n161), .Y(n162) );
  OAI22XL U622 ( .A0(n312), .A1(n221), .B0(n514), .B1(n225), .Y(n390) );
  AOI21X1 U623 ( .A0(n312), .A1(n226), .B0(n227), .Y(n225) );
  NAND4X1 U624 ( .A(n211), .B(n121), .C(n535), .D(n47), .Y(n226) );
  OAI22XL U625 ( .A0(n318), .A1(n105), .B0(n502), .B1(n116), .Y(n360) );
  AOI222XL U626 ( .A0(n117), .A1(n109), .B0(N185), .B1(n110), .C0(n508), .C1(
        n112), .Y(n116) );
  OAI22XL U627 ( .A0(n322), .A1(n156), .B0(n504), .B1(n163), .Y(n372) );
  AOI222XL U628 ( .A0(n117), .A1(n159), .B0(N185), .B1(n160), .C0(n508), .C1(
        n161), .Y(n163) );
  OAI22XL U629 ( .A0(n282), .A1(n156), .B0(n504), .B1(n158), .Y(n370) );
  AOI222XL U630 ( .A0(n108), .A1(n159), .B0(N183), .B1(n160), .C0(n506), .C1(
        n161), .Y(n158) );
  OAI22XL U631 ( .A0(n514), .A1(n223), .B0(n310), .B1(n238), .Y(n395) );
  NOR2X1 U632 ( .A(n514), .B(n196), .Y(n238) );
  NAND2X1 U633 ( .A(n334), .B(n335), .Y(n145) );
  OAI22XL U634 ( .A0(n328), .A1(n173), .B0(n505), .B1(n182), .Y(n378) );
  AOI221XL U635 ( .A0(n508), .A1(n176), .B0(n177), .B1(N185), .C0(n117), .Y(
        n182) );
  OAI22XL U636 ( .A0(n327), .A1(n173), .B0(n505), .B1(n180), .Y(n377) );
  AOI221XL U637 ( .A0(n507), .A1(n176), .B0(n177), .B1(n441), .C0(n114), .Y(
        n180) );
  OAI22XL U638 ( .A0(n326), .A1(n173), .B0(n505), .B1(n175), .Y(n376) );
  AOI221XL U639 ( .A0(n506), .A1(n176), .B0(n177), .B1(N183), .C0(n108), .Y(
        n175) );
  OAI22XL U640 ( .A0(n518), .A1(n81), .B0(n82), .B1(n294), .Y(n343) );
  AOI222XL U641 ( .A0(n537), .A1(\buff[7][2] ), .B0(n86), .B1(n294), .C0(N180), 
        .C1(n79), .Y(n81) );
  OA21XL U642 ( .A0(n331), .A1(n83), .B0(n84), .Y(n82) );
  AOI2BB1X1 U643 ( .A0N(n315), .A1N(n83), .B0(n518), .Y(n234) );
  CLKINVX1 U644 ( .A(n334), .Y(n542) );
  NAND2X1 U645 ( .A(n334), .B(N156), .Y(n135) );
  OAI21XL U646 ( .A0(n311), .A1(n221), .B0(n222), .Y(n389) );
  OAI2BB1X1 U647 ( .A0N(n223), .A1N(n189), .B0(n221), .Y(n222) );
  OA21XL U648 ( .A0(n332), .A1(n83), .B0(n89), .Y(n84) );
  OAI211X1 U649 ( .A0(n290), .A1(n250), .B0(n256), .C0(n519), .Y(n241) );
  OA22X1 U650 ( .A0(n130), .A1(n286), .B0(n288), .B1(n109), .Y(n256) );
  CLKINVX1 U651 ( .A(n258), .Y(n519) );
  OAI221XL U652 ( .A0(n140), .A1(n284), .B0(n149), .B1(n282), .C0(n259), .Y(
        n258) );
  OAI211X1 U653 ( .A0(n289), .A1(n250), .B0(n252), .C0(n520), .Y(n251) );
  OA22X1 U654 ( .A0(n130), .A1(n285), .B0(n287), .B1(n109), .Y(n252) );
  CLKINVX1 U655 ( .A(n254), .Y(n520) );
  OAI221XL U656 ( .A0(n140), .A1(n283), .B0(n149), .B1(n281), .C0(n255), .Y(
        n254) );
  NAND3X1 U657 ( .A(n231), .B(n42), .C(n236), .Y(n394) );
  AOI2BB2X1 U658 ( .B0(n237), .B1(W[2]), .A0N(n535), .A1N(n310), .Y(n236) );
  OAI21XL U659 ( .A0(n314), .A1(n83), .B0(n234), .Y(n237) );
  OA22X1 U660 ( .A0(n323), .A1(n159), .B0(n326), .B1(n168), .Y(n259) );
  OA22X1 U661 ( .A0(n324), .A1(n159), .B0(n327), .B1(n168), .Y(n255) );
  CLKBUFX3 U662 ( .A(N184), .Y(n441) );
  MXI2X1 U663 ( .A(n449), .B(n450), .S0(N158), .Y(N184) );
  MXI4X1 U664 ( .A(\buff[0][1] ), .B(\buff[1][1] ), .C(\buff[2][1] ), .D(
        \buff[3][1] ), .S0(N156), .S1(N157), .Y(n449) );
  MXI4X1 U665 ( .A(\buff[4][1] ), .B(\buff[5][1] ), .C(\buff[6][1] ), .D(
        \buff[7][1] ), .S0(N156), .S1(N157), .Y(n450) );
  AO22X1 U666 ( .A0(state[0]), .A1(n516), .B0(n213), .B1(n214), .Y(n387) );
  AO21X1 U667 ( .A0(n215), .A1(n198), .B0(n183), .Y(n213) );
  NAND2X2 U668 ( .A(n317), .B(n316), .Y(n83) );
  NOR2X2 U669 ( .A(n400), .B(n316), .Y(n79) );
  OAI211X1 U670 ( .A0(n315), .A1(n89), .B0(n231), .C0(n235), .Y(n393) );
  AOI2BB2X1 U671 ( .B0(n315), .B1(n538), .A0N(n535), .A1N(n312), .Y(n235) );
  OAI22XL U672 ( .A0(n399), .A1(n214), .B0(n516), .B1(n217), .Y(n388) );
  AOI2BB1X1 U673 ( .A0N(state[1]), .A1N(n530), .B0(n183), .Y(n217) );
  CLKINVX1 U674 ( .A(n46), .Y(n521) );
  OAI32XL U675 ( .A0(Valid), .A1(n316), .A2(n317), .B0(n47), .B1(n522), .Y(n46) );
  OAI2BB2XL U676 ( .B0(n332), .B1(n89), .A0N(n89), .A1N(n93), .Y(n345) );
  OAI221XL U677 ( .A0(n91), .A1(n291), .B0(n398), .B1(n535), .C0(n88), .Y(n93)
         );
  NAND2X1 U678 ( .A(N251), .B(n181), .Y(n179) );
  MXI2X1 U679 ( .A(n455), .B(n456), .S0(N161), .Y(N251) );
  MXI4X1 U680 ( .A(\buff[4][2] ), .B(\buff[5][2] ), .C(\buff[6][2] ), .D(
        \buff[7][2] ), .S0(N159), .S1(N160), .Y(n456) );
  MXI4X1 U681 ( .A(\buff[0][2] ), .B(\buff[1][2] ), .C(\buff[2][2] ), .D(
        \buff[3][2] ), .S0(N159), .S1(N160), .Y(n455) );
  NAND2X1 U682 ( .A(N253), .B(n181), .Y(n103) );
  MXI2X1 U683 ( .A(n451), .B(n452), .S0(N161), .Y(N253) );
  MXI4X1 U684 ( .A(\buff[4][0] ), .B(\buff[5][0] ), .C(\buff[6][0] ), .D(
        \buff[7][0] ), .S0(N159), .S1(N160), .Y(n452) );
  MXI4X1 U685 ( .A(\buff[0][0] ), .B(\buff[1][0] ), .C(\buff[2][0] ), .D(
        \buff[3][0] ), .S0(N159), .S1(N160), .Y(n451) );
  NAND2X1 U686 ( .A(N252), .B(n181), .Y(n98) );
  MXI2X1 U687 ( .A(n453), .B(n454), .S0(N161), .Y(N252) );
  MXI4X1 U688 ( .A(\buff[4][1] ), .B(\buff[5][1] ), .C(\buff[6][1] ), .D(
        \buff[7][1] ), .S0(N159), .S1(N160), .Y(n454) );
  MXI4X1 U689 ( .A(\buff[0][1] ), .B(\buff[1][1] ), .C(\buff[2][1] ), .D(
        \buff[3][1] ), .S0(N159), .S1(N160), .Y(n453) );
  OAI2BB2XL U690 ( .B0(n309), .B1(n228), .A0N(n534), .A1N(n228), .Y(n391) );
  OAI31XL U691 ( .A0(W[2]), .A1(n535), .A2(n230), .B0(n41), .Y(n228) );
  OAI2BB2XL U692 ( .B0(n331), .B1(n84), .A0N(n89), .A1N(n90), .Y(n344) );
  OAI222XL U693 ( .A0(n91), .A1(n292), .B0(J[1]), .B1(n88), .C0(n524), .C1(
        n535), .Y(n90) );
  NAND3BX1 U694 ( .AN(n230), .B(n538), .C(n313), .Y(n42) );
  NAND2X1 U695 ( .A(n332), .B(n538), .Y(n88) );
  NAND2X1 U696 ( .A(n314), .B(n315), .Y(n230) );
  OA21XL U697 ( .A0(n311), .A1(n312), .B0(n196), .Y(n189) );
  CLKINVX1 U698 ( .A(\val[2] ), .Y(n539) );
  OAI22XL U699 ( .A0(sum[1]), .A1(n457), .B0(n457), .B1(n408), .Y(n459) );
  NAND2X1 U700 ( .A(sum[7]), .B(n480), .Y(n471) );
  NAND2X1 U701 ( .A(sum[6]), .B(n479), .Y(n466) );
  NOR3BXL U702 ( .AN(n466), .B(n460), .C(n467), .Y(n458) );
  NAND3X1 U703 ( .A(n459), .B(n471), .C(n458), .Y(n478) );
  NAND2X1 U704 ( .A(sum[9]), .B(n401), .Y(n474) );
  NAND2X1 U705 ( .A(sum[2]), .B(n430), .Y(n473) );
  OAI211X1 U706 ( .A0(n462), .A1(n485), .B0(n461), .C0(n473), .Y(n463) );
  OAI221XL U707 ( .A0(sum[2]), .A1(n430), .B0(sum[3]), .B1(n423), .C0(n463), 
        .Y(n464) );
  NOR4X1 U708 ( .A(n478), .B(n477), .C(n476), .D(n475), .Y(N452) );
endmodule

