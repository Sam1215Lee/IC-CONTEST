
module LCD_CTRL_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
endmodule


module LCD_CTRL ( clk, reset, datain, cmd, cmd_valid, dataout, output_valid, 
        busy );
  input [7:0] datain;
  input [2:0] cmd;
  output [7:0] dataout;
  input clk, reset, cmd_valid;
  output output_valid, busy;
  wire   next_state, N966, N971, N972, N973, N981, N982, N983, N984, N987,
         N988, N999, N1000, N1001, N1002, N1003, \img_buff[0][7] ,
         \img_buff[0][6] , \img_buff[0][5] , \img_buff[0][4] ,
         \img_buff[0][3] , \img_buff[0][2] , \img_buff[0][1] ,
         \img_buff[0][0] , \img_buff[2][7] , \img_buff[2][6] ,
         \img_buff[2][5] , \img_buff[2][4] , \img_buff[2][3] ,
         \img_buff[2][2] , \img_buff[2][1] , \img_buff[2][0] ,
         \img_buff[4][7] , \img_buff[4][6] , \img_buff[4][5] ,
         \img_buff[4][4] , \img_buff[4][3] , \img_buff[4][2] ,
         \img_buff[4][1] , \img_buff[4][0] , \img_buff[5][7] ,
         \img_buff[5][6] , \img_buff[5][5] , \img_buff[5][4] ,
         \img_buff[5][3] , \img_buff[5][2] , \img_buff[5][1] ,
         \img_buff[5][0] , \img_buff[6][7] , \img_buff[6][6] ,
         \img_buff[6][5] , \img_buff[6][4] , \img_buff[6][3] ,
         \img_buff[6][2] , \img_buff[6][1] , \img_buff[6][0] ,
         \img_buff[7][7] , \img_buff[7][6] , \img_buff[7][5] ,
         \img_buff[7][4] , \img_buff[7][3] , \img_buff[7][2] ,
         \img_buff[7][1] , \img_buff[7][0] , \img_buff[8][7] ,
         \img_buff[8][6] , \img_buff[8][5] , \img_buff[8][4] ,
         \img_buff[8][3] , \img_buff[8][2] , \img_buff[8][1] ,
         \img_buff[8][0] , \img_buff[11][7] , \img_buff[11][6] ,
         \img_buff[11][5] , \img_buff[11][4] , \img_buff[11][3] ,
         \img_buff[11][2] , \img_buff[11][1] , \img_buff[11][0] ,
         \img_buff[12][7] , \img_buff[12][6] , \img_buff[12][5] ,
         \img_buff[12][4] , \img_buff[12][3] , \img_buff[12][2] ,
         \img_buff[12][1] , \img_buff[12][0] , \img_buff[13][7] ,
         \img_buff[13][6] , \img_buff[13][5] , \img_buff[13][4] ,
         \img_buff[13][3] , \img_buff[13][2] , \img_buff[13][1] ,
         \img_buff[13][0] , \img_buff[14][7] , \img_buff[14][6] ,
         \img_buff[14][5] , \img_buff[14][4] , \img_buff[14][3] ,
         \img_buff[14][2] , \img_buff[14][1] , \img_buff[14][0] ,
         \img_buff[15][7] , \img_buff[15][6] , \img_buff[15][5] ,
         \img_buff[15][4] , \img_buff[15][3] , \img_buff[15][2] ,
         \img_buff[15][1] , \img_buff[15][0] , \img_buff[16][7] ,
         \img_buff[16][6] , \img_buff[16][5] , \img_buff[16][4] ,
         \img_buff[16][3] , \img_buff[16][2] , \img_buff[16][1] ,
         \img_buff[16][0] , \img_buff[17][7] , \img_buff[17][6] ,
         \img_buff[17][5] , \img_buff[17][4] , \img_buff[17][3] ,
         \img_buff[17][2] , \img_buff[17][1] , \img_buff[17][0] ,
         \img_buff[20][7] , \img_buff[20][6] , \img_buff[20][5] ,
         \img_buff[20][4] , \img_buff[20][3] , \img_buff[20][2] ,
         \img_buff[20][1] , \img_buff[20][0] , \img_buff[22][7] ,
         \img_buff[22][6] , \img_buff[22][5] , \img_buff[22][4] ,
         \img_buff[22][3] , \img_buff[22][2] , \img_buff[22][1] ,
         \img_buff[22][0] , \img_buff[23][7] , \img_buff[23][6] ,
         \img_buff[23][5] , \img_buff[23][4] , \img_buff[23][3] ,
         \img_buff[23][2] , \img_buff[23][1] , \img_buff[23][0] ,
         \img_buff[27][7] , \img_buff[27][6] , \img_buff[27][5] ,
         \img_buff[27][4] , \img_buff[27][3] , \img_buff[27][2] ,
         \img_buff[27][1] , \img_buff[27][0] , \img_buff[28][7] ,
         \img_buff[28][6] , \img_buff[28][5] , \img_buff[28][4] ,
         \img_buff[28][3] , \img_buff[28][2] , \img_buff[28][1] ,
         \img_buff[28][0] , \img_buff[29][7] , \img_buff[29][6] ,
         \img_buff[29][5] , \img_buff[29][4] , \img_buff[29][3] ,
         \img_buff[29][2] , \img_buff[29][1] , \img_buff[29][0] ,
         \img_buff[30][7] , \img_buff[30][6] , \img_buff[30][5] ,
         \img_buff[30][4] , \img_buff[30][3] , \img_buff[30][2] ,
         \img_buff[30][1] , \img_buff[30][0] , \img_buff[33][7] ,
         \img_buff[33][6] , \img_buff[33][5] , \img_buff[33][4] ,
         \img_buff[33][3] , \img_buff[33][2] , \img_buff[33][1] ,
         \img_buff[33][0] , \img_buff[34][7] , \img_buff[34][6] ,
         \img_buff[34][5] , \img_buff[34][4] , \img_buff[34][3] ,
         \img_buff[34][2] , \img_buff[34][1] , \img_buff[34][0] ,
         \img_buff[35][7] , \img_buff[35][6] , \img_buff[35][5] ,
         \img_buff[35][4] , \img_buff[35][3] , \img_buff[35][2] ,
         \img_buff[35][1] , \img_buff[35][0] , \img_buff[38][7] ,
         \img_buff[38][6] , \img_buff[38][5] , \img_buff[38][4] ,
         \img_buff[38][3] , \img_buff[38][2] , \img_buff[38][1] ,
         \img_buff[38][0] , \img_buff[39][7] , \img_buff[39][6] ,
         \img_buff[39][5] , \img_buff[39][4] , \img_buff[39][3] ,
         \img_buff[39][2] , \img_buff[39][1] , \img_buff[39][0] ,
         \img_buff[40][7] , \img_buff[40][6] , \img_buff[40][5] ,
         \img_buff[40][4] , \img_buff[40][3] , \img_buff[40][2] ,
         \img_buff[40][1] , \img_buff[40][0] , \img_buff[41][7] ,
         \img_buff[41][6] , \img_buff[41][5] , \img_buff[41][4] ,
         \img_buff[41][3] , \img_buff[41][2] , \img_buff[41][1] ,
         \img_buff[41][0] , \img_buff[42][7] , \img_buff[42][6] ,
         \img_buff[42][5] , \img_buff[42][4] , \img_buff[42][3] ,
         \img_buff[42][2] , \img_buff[42][1] , \img_buff[42][0] ,
         \img_buff[43][7] , \img_buff[43][6] , \img_buff[43][5] ,
         \img_buff[43][4] , \img_buff[43][3] , \img_buff[43][2] ,
         \img_buff[43][1] , \img_buff[43][0] , \img_buff[44][7] ,
         \img_buff[44][6] , \img_buff[44][5] , \img_buff[44][4] ,
         \img_buff[44][3] , \img_buff[44][2] , \img_buff[44][1] ,
         \img_buff[44][0] , \img_buff[47][7] , \img_buff[47][6] ,
         \img_buff[47][5] , \img_buff[47][4] , \img_buff[47][3] ,
         \img_buff[47][2] , \img_buff[47][1] , \img_buff[47][0] ,
         \img_buff[49][7] , \img_buff[49][6] , \img_buff[49][5] ,
         \img_buff[49][4] , \img_buff[49][3] , \img_buff[49][2] ,
         \img_buff[49][1] , \img_buff[49][0] , \img_buff[50][7] ,
         \img_buff[50][6] , \img_buff[50][5] , \img_buff[50][4] ,
         \img_buff[50][3] , \img_buff[50][2] , \img_buff[50][1] ,
         \img_buff[50][0] , \img_buff[54][7] , \img_buff[54][6] ,
         \img_buff[54][5] , \img_buff[54][4] , \img_buff[54][3] ,
         \img_buff[54][2] , \img_buff[54][1] , \img_buff[54][0] ,
         \img_buff[55][7] , \img_buff[55][6] , \img_buff[55][5] ,
         \img_buff[55][4] , \img_buff[55][3] , \img_buff[55][2] ,
         \img_buff[55][1] , \img_buff[55][0] , \img_buff[56][7] ,
         \img_buff[56][6] , \img_buff[56][5] , \img_buff[56][4] ,
         \img_buff[56][3] , \img_buff[56][2] , \img_buff[56][1] ,
         \img_buff[56][0] , \img_buff[57][7] , \img_buff[57][6] ,
         \img_buff[57][5] , \img_buff[57][4] , \img_buff[57][3] ,
         \img_buff[57][2] , \img_buff[57][1] , \img_buff[57][0] ,
         \img_buff[60][7] , \img_buff[60][6] , \img_buff[60][5] ,
         \img_buff[60][4] , \img_buff[60][3] , \img_buff[60][2] ,
         \img_buff[60][1] , \img_buff[60][0] , \img_buff[61][7] ,
         \img_buff[61][6] , \img_buff[61][5] , \img_buff[61][4] ,
         \img_buff[61][3] , \img_buff[61][2] , \img_buff[61][1] ,
         \img_buff[61][0] , \img_buff[62][7] , \img_buff[62][6] ,
         \img_buff[62][5] , \img_buff[62][4] , \img_buff[62][3] ,
         \img_buff[62][2] , \img_buff[62][1] , \img_buff[62][0] ,
         \img_buff[63][7] , \img_buff[63][6] , \img_buff[63][5] ,
         \img_buff[63][4] , \img_buff[63][3] , \img_buff[63][2] ,
         \img_buff[63][1] , \img_buff[63][0] , \img_buff[64][7] ,
         \img_buff[64][6] , \img_buff[64][5] , \img_buff[64][4] ,
         \img_buff[64][3] , \img_buff[64][2] , \img_buff[64][1] ,
         \img_buff[64][0] , \img_buff[67][7] , \img_buff[67][6] ,
         \img_buff[67][5] , \img_buff[67][4] , \img_buff[67][3] ,
         \img_buff[67][2] , \img_buff[67][1] , \img_buff[67][0] ,
         \img_buff[68][7] , \img_buff[68][6] , \img_buff[68][5] ,
         \img_buff[68][4] , \img_buff[68][3] , \img_buff[68][2] ,
         \img_buff[68][1] , \img_buff[68][0] , \img_buff[69][7] ,
         \img_buff[69][6] , \img_buff[69][5] , \img_buff[69][4] ,
         \img_buff[69][3] , \img_buff[69][2] , \img_buff[69][1] ,
         \img_buff[69][0] , \img_buff[72][7] , \img_buff[72][6] ,
         \img_buff[72][5] , \img_buff[72][4] , \img_buff[72][3] ,
         \img_buff[72][2] , \img_buff[72][1] , \img_buff[72][0] ,
         \img_buff[73][7] , \img_buff[73][6] , \img_buff[73][5] ,
         \img_buff[73][4] , \img_buff[73][3] , \img_buff[73][2] ,
         \img_buff[73][1] , \img_buff[73][0] , \img_buff[74][7] ,
         \img_buff[74][6] , \img_buff[74][5] , \img_buff[74][4] ,
         \img_buff[74][3] , \img_buff[74][2] , \img_buff[74][1] ,
         \img_buff[74][0] , \img_buff[76][7] , \img_buff[76][6] ,
         \img_buff[76][5] , \img_buff[76][4] , \img_buff[76][3] ,
         \img_buff[76][2] , \img_buff[76][1] , \img_buff[76][0] ,
         \img_buff[79][7] , \img_buff[79][6] , \img_buff[79][5] ,
         \img_buff[79][4] , \img_buff[79][3] , \img_buff[79][2] ,
         \img_buff[79][1] , \img_buff[79][0] , \img_buff[81][7] ,
         \img_buff[81][6] , \img_buff[81][5] , \img_buff[81][4] ,
         \img_buff[81][3] , \img_buff[81][2] , \img_buff[81][1] ,
         \img_buff[81][0] , \img_buff[82][7] , \img_buff[82][6] ,
         \img_buff[82][5] , \img_buff[82][4] , \img_buff[82][3] ,
         \img_buff[82][2] , \img_buff[82][1] , \img_buff[82][0] ,
         \img_buff[83][7] , \img_buff[83][6] , \img_buff[83][5] ,
         \img_buff[83][4] , \img_buff[83][3] , \img_buff[83][2] ,
         \img_buff[83][1] , \img_buff[83][0] , \img_buff[84][7] ,
         \img_buff[84][6] , \img_buff[84][5] , \img_buff[84][4] ,
         \img_buff[84][3] , \img_buff[84][2] , \img_buff[84][1] ,
         \img_buff[84][0] , \img_buff[87][7] , \img_buff[87][6] ,
         \img_buff[87][5] , \img_buff[87][4] , \img_buff[87][3] ,
         \img_buff[87][2] , \img_buff[87][1] , \img_buff[87][0] ,
         \img_buff[88][7] , \img_buff[88][6] , \img_buff[88][5] ,
         \img_buff[88][4] , \img_buff[88][3] , \img_buff[88][2] ,
         \img_buff[88][1] , \img_buff[88][0] , \img_buff[89][7] ,
         \img_buff[89][6] , \img_buff[89][5] , \img_buff[89][4] ,
         \img_buff[89][3] , \img_buff[89][2] , \img_buff[89][1] ,
         \img_buff[89][0] , \img_buff[94][7] , \img_buff[94][6] ,
         \img_buff[94][5] , \img_buff[94][4] , \img_buff[94][3] ,
         \img_buff[94][2] , \img_buff[94][1] , \img_buff[94][0] ,
         \img_buff[95][7] , \img_buff[95][6] , \img_buff[95][5] ,
         \img_buff[95][4] , \img_buff[95][3] , \img_buff[95][2] ,
         \img_buff[95][1] , \img_buff[95][0] , \img_buff[96][7] ,
         \img_buff[96][6] , \img_buff[96][5] , \img_buff[96][4] ,
         \img_buff[96][3] , \img_buff[96][2] , \img_buff[96][1] ,
         \img_buff[96][0] , \img_buff[97][7] , \img_buff[97][6] ,
         \img_buff[97][5] , \img_buff[97][4] , \img_buff[97][3] ,
         \img_buff[97][2] , \img_buff[97][1] , \img_buff[97][0] ,
         \img_buff[98][7] , \img_buff[98][6] , \img_buff[98][5] ,
         \img_buff[98][4] , \img_buff[98][3] , \img_buff[98][2] ,
         \img_buff[98][1] , \img_buff[98][0] , \img_buff[101][7] ,
         \img_buff[101][6] , \img_buff[101][5] , \img_buff[101][4] ,
         \img_buff[101][3] , \img_buff[101][2] , \img_buff[101][1] ,
         \img_buff[101][0] , \img_buff[102][7] , \img_buff[102][6] ,
         \img_buff[102][5] , \img_buff[102][4] , \img_buff[102][3] ,
         \img_buff[102][2] , \img_buff[102][1] , \img_buff[102][0] ,
         \img_buff[103][7] , \img_buff[103][6] , \img_buff[103][5] ,
         \img_buff[103][4] , \img_buff[103][3] , \img_buff[103][2] ,
         \img_buff[103][1] , \img_buff[103][0] , \img_buff[107][7] ,
         \img_buff[107][6] , \img_buff[107][5] , \img_buff[107][4] ,
         \img_buff[107][3] , \img_buff[107][2] , \img_buff[107][1] ,
         \img_buff[107][0] , N1160, N1161, N1162, N1163, N1164, N1165, N1166,
         N1167, \U3/U10/Z_1 , \U3/U10/Z_2 , \U3/U10/Z_3 , \U3/U11/Z_0 ,
         \U3/U11/Z_1 , \U3/U11/Z_2 , \U3/U11/Z_3 , \U3/U12/Z_4 , \U3/U12/Z_5 ,
         \U3/U12/Z_6 , \U3/U13/Z_2 , \U3/U13/Z_3 , \U3/U15/Z_3 , \U3/U15/Z_4 ,
         \U3/U15/Z_5 , \U3/U15/Z_6 , \U3/U16/Z_4 , \U3/U16/Z_5 , \U3/U16/Z_6 ,
         n205, n216, n217, n218, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n408, n409, n410, n411, n412, n413,
         n414, n415, n424, n425, n426, n429, n430, n431, n432, n1236, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, \r481/carry[6] ,
         \r481/carry[5] , \r481/carry[4] , \r481/carry[3] , \r594/carry[6] ,
         \r594/carry[5] , \r594/carry[4] , \r596/carry[6] , \r596/carry[5] ,
         \r596/carry[4] , \r596/carry[3] , \r596/carry[2] , \r596/carry[1] ,
         \r597/carry[4] , \r597/carry[3] , \r597/carry[2] , \r597/carry[1] ,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418;
  wire   [7:0] img_counter;
  wire   [6:0] out_pos;

  LCD_CTRL_DW01_inc_0 r452 ( .A(img_counter), .SUM({N1167, N1166, N1165, N1164, 
        N1163, N1162, N1161, N1160}) );
  EDFFX1 mode_reg ( .D(n2418), .E(n1236), .CK(clk), .Q(n1290), .QN(n432) );
  DFFRXL \W_reg[1]  ( .D(n1280), .CK(clk), .RN(n2309), .QN(n430) );
  DFFRXL cur_state_reg ( .D(next_state), .CK(clk), .RN(n2309), .Q(n1284), .QN(
        n205) );
  DFFRXL \L_reg[3]  ( .D(n1262), .CK(clk), .RN(n2309), .QN(n424) );
  EDFFX1 \img_buff_reg[1][7]  ( .D(datain[7]), .E(n2416), .CK(clk), .QN(n2287)
         );
  EDFFX1 \img_buff_reg[1][6]  ( .D(datain[6]), .E(n2416), .CK(clk), .QN(n2253)
         );
  EDFFX1 \img_buff_reg[1][5]  ( .D(datain[5]), .E(n2416), .CK(clk), .QN(n2219)
         );
  EDFFX1 \img_buff_reg[1][4]  ( .D(datain[4]), .E(n2416), .CK(clk), .QN(n2185)
         );
  EDFFX1 \img_buff_reg[1][3]  ( .D(datain[3]), .E(n2416), .CK(clk), .QN(n2151)
         );
  EDFFX1 \img_buff_reg[1][2]  ( .D(datain[2]), .E(n2416), .CK(clk), .QN(n2117)
         );
  EDFFX1 \img_buff_reg[1][1]  ( .D(datain[1]), .E(n2416), .CK(clk), .QN(n2083)
         );
  EDFFX1 \img_buff_reg[1][0]  ( .D(datain[0]), .E(n2416), .CK(clk), .QN(n2049)
         );
  EDFFX1 \img_buff_reg[3][7]  ( .D(datain[7]), .E(n2414), .CK(clk), .QN(n2286)
         );
  EDFFX1 \img_buff_reg[3][6]  ( .D(datain[6]), .E(n2414), .CK(clk), .QN(n2252)
         );
  EDFFX1 \img_buff_reg[3][5]  ( .D(datain[5]), .E(n2414), .CK(clk), .QN(n2218)
         );
  EDFFX1 \img_buff_reg[3][4]  ( .D(datain[4]), .E(n2414), .CK(clk), .QN(n2184)
         );
  EDFFX1 \img_buff_reg[3][3]  ( .D(datain[3]), .E(n2414), .CK(clk), .QN(n2150)
         );
  EDFFX1 \img_buff_reg[3][2]  ( .D(datain[2]), .E(n2414), .CK(clk), .QN(n2116)
         );
  EDFFX1 \img_buff_reg[3][1]  ( .D(datain[1]), .E(n2414), .CK(clk), .QN(n2082)
         );
  EDFFX1 \img_buff_reg[3][0]  ( .D(datain[0]), .E(n2414), .CK(clk), .QN(n2048)
         );
  EDFFX1 \img_buff_reg[9][7]  ( .D(datain[7]), .E(n2408), .CK(clk), .QN(n232)
         );
  EDFFX1 \img_buff_reg[9][6]  ( .D(datain[6]), .E(n2408), .CK(clk), .QN(n233)
         );
  EDFFX1 \img_buff_reg[9][5]  ( .D(datain[5]), .E(n2408), .CK(clk), .QN(n234)
         );
  EDFFX1 \img_buff_reg[9][4]  ( .D(datain[4]), .E(n2408), .CK(clk), .QN(n235)
         );
  EDFFX1 \img_buff_reg[9][3]  ( .D(datain[3]), .E(n2408), .CK(clk), .QN(n236)
         );
  EDFFX1 \img_buff_reg[9][2]  ( .D(datain[2]), .E(n2408), .CK(clk), .QN(n237)
         );
  EDFFX1 \img_buff_reg[9][1]  ( .D(datain[1]), .E(n2408), .CK(clk), .QN(n238)
         );
  EDFFX1 \img_buff_reg[9][0]  ( .D(datain[0]), .E(n2408), .CK(clk), .QN(n239)
         );
  EDFFX1 \img_buff_reg[10][7]  ( .D(datain[7]), .E(n2407), .CK(clk), .QN(n240)
         );
  EDFFX1 \img_buff_reg[10][6]  ( .D(datain[6]), .E(n2407), .CK(clk), .QN(n241)
         );
  EDFFX1 \img_buff_reg[10][5]  ( .D(datain[5]), .E(n2407), .CK(clk), .QN(n242)
         );
  EDFFX1 \img_buff_reg[10][4]  ( .D(datain[4]), .E(n2407), .CK(clk), .QN(n243)
         );
  EDFFX1 \img_buff_reg[10][3]  ( .D(datain[3]), .E(n2407), .CK(clk), .QN(n244)
         );
  EDFFX1 \img_buff_reg[10][2]  ( .D(datain[2]), .E(n2407), .CK(clk), .QN(n245)
         );
  EDFFX1 \img_buff_reg[10][1]  ( .D(datain[1]), .E(n2407), .CK(clk), .QN(n246)
         );
  EDFFX1 \img_buff_reg[10][0]  ( .D(datain[0]), .E(n2407), .CK(clk), .QN(n247)
         );
  EDFFX1 \img_buff_reg[21][4]  ( .D(datain[4]), .E(n2396), .CK(clk), .QN(n2189) );
  EDFFX1 \img_buff_reg[21][3]  ( .D(datain[3]), .E(n2396), .CK(clk), .QN(n2155) );
  EDFFX1 \img_buff_reg[21][2]  ( .D(datain[2]), .E(n2396), .CK(clk), .QN(n2121) );
  EDFFX1 \img_buff_reg[21][1]  ( .D(datain[1]), .E(n2396), .CK(clk), .QN(n2087) );
  EDFFX1 \img_buff_reg[21][0]  ( .D(datain[0]), .E(n2396), .CK(clk), .QN(n2053) );
  EDFFX1 \img_buff_reg[21][7]  ( .D(datain[7]), .E(n2396), .CK(clk), .QN(n2291) );
  EDFFX1 \img_buff_reg[21][6]  ( .D(datain[6]), .E(n2396), .CK(clk), .QN(n2257) );
  EDFFX1 \img_buff_reg[21][5]  ( .D(datain[5]), .E(n2396), .CK(clk), .QN(n2223) );
  EDFFX1 \img_buff_reg[24][7]  ( .D(datain[7]), .E(n2393), .CK(clk), .QN(n2288) );
  EDFFX1 \img_buff_reg[24][6]  ( .D(datain[6]), .E(n2393), .CK(clk), .QN(n2254) );
  EDFFX1 \img_buff_reg[24][5]  ( .D(datain[5]), .E(n2393), .CK(clk), .QN(n2220) );
  EDFFX1 \img_buff_reg[24][4]  ( .D(datain[4]), .E(n2393), .CK(clk), .QN(n2186) );
  EDFFX1 \img_buff_reg[24][3]  ( .D(datain[3]), .E(n2393), .CK(clk), .QN(n2152) );
  EDFFX1 \img_buff_reg[24][2]  ( .D(datain[2]), .E(n2393), .CK(clk), .QN(n2118) );
  EDFFX1 \img_buff_reg[24][1]  ( .D(datain[1]), .E(n2393), .CK(clk), .QN(n2084) );
  EDFFX1 \img_buff_reg[24][0]  ( .D(datain[0]), .E(n2393), .CK(clk), .QN(n2050) );
  EDFFX1 \img_buff_reg[31][7]  ( .D(datain[7]), .E(n2386), .CK(clk), .QN(n2294) );
  EDFFX1 \img_buff_reg[31][6]  ( .D(datain[6]), .E(n2386), .CK(clk), .QN(n2260) );
  EDFFX1 \img_buff_reg[31][5]  ( .D(datain[5]), .E(n2386), .CK(clk), .QN(n2226) );
  EDFFX1 \img_buff_reg[31][4]  ( .D(datain[4]), .E(n2386), .CK(clk), .QN(n2192) );
  EDFFX1 \img_buff_reg[31][3]  ( .D(datain[3]), .E(n2386), .CK(clk), .QN(n2158) );
  EDFFX1 \img_buff_reg[31][2]  ( .D(datain[2]), .E(n2386), .CK(clk), .QN(n2124) );
  EDFFX1 \img_buff_reg[31][1]  ( .D(datain[1]), .E(n2386), .CK(clk), .QN(n2090) );
  EDFFX1 \img_buff_reg[31][0]  ( .D(datain[0]), .E(n2386), .CK(clk), .QN(n2056) );
  EDFFX1 \img_buff_reg[48][7]  ( .D(datain[7]), .E(n2369), .CK(clk), .QN(n2299) );
  EDFFX1 \img_buff_reg[48][6]  ( .D(datain[6]), .E(n2369), .CK(clk), .QN(n2265) );
  EDFFX1 \img_buff_reg[48][5]  ( .D(datain[5]), .E(n2369), .CK(clk), .QN(n2231) );
  EDFFX1 \img_buff_reg[48][4]  ( .D(datain[4]), .E(n2369), .CK(clk), .QN(n2197) );
  EDFFX1 \img_buff_reg[48][3]  ( .D(datain[3]), .E(n2369), .CK(clk), .QN(n2163) );
  EDFFX1 \img_buff_reg[48][2]  ( .D(datain[2]), .E(n2369), .CK(clk), .QN(n2129) );
  EDFFX1 \img_buff_reg[48][1]  ( .D(datain[1]), .E(n2369), .CK(clk), .QN(n2095) );
  EDFFX1 \img_buff_reg[48][0]  ( .D(datain[0]), .E(n2369), .CK(clk), .QN(n2061) );
  EDFFX1 \img_buff_reg[51][7]  ( .D(datain[7]), .E(n2366), .CK(clk), .QN(n2296) );
  EDFFX1 \img_buff_reg[51][6]  ( .D(datain[6]), .E(n2366), .CK(clk), .QN(n2262) );
  EDFFX1 \img_buff_reg[51][5]  ( .D(datain[5]), .E(n2366), .CK(clk), .QN(n2228) );
  EDFFX1 \img_buff_reg[51][4]  ( .D(datain[4]), .E(n2366), .CK(clk), .QN(n2194) );
  EDFFX1 \img_buff_reg[51][3]  ( .D(datain[3]), .E(n2366), .CK(clk), .QN(n2160) );
  EDFFX1 \img_buff_reg[51][2]  ( .D(datain[2]), .E(n2366), .CK(clk), .QN(n2126) );
  EDFFX1 \img_buff_reg[51][1]  ( .D(datain[1]), .E(n2366), .CK(clk), .QN(n2092) );
  EDFFX1 \img_buff_reg[51][0]  ( .D(datain[0]), .E(n2366), .CK(clk), .QN(n2058) );
  EDFFX1 \img_buff_reg[58][3]  ( .D(datain[3]), .E(n2359), .CK(clk), .QN(n2132) );
  EDFFX1 \img_buff_reg[58][2]  ( .D(datain[2]), .E(n2359), .CK(clk), .QN(n2098) );
  EDFFX1 \img_buff_reg[58][1]  ( .D(datain[1]), .E(n2359), .CK(clk), .QN(n2064) );
  EDFFX1 \img_buff_reg[58][0]  ( .D(datain[0]), .E(n2359), .CK(clk), .QN(n2030) );
  EDFFX1 \img_buff_reg[58][7]  ( .D(datain[7]), .E(n2359), .CK(clk), .QN(n2268) );
  EDFFX1 \img_buff_reg[58][6]  ( .D(datain[6]), .E(n2359), .CK(clk), .QN(n2234) );
  EDFFX1 \img_buff_reg[58][5]  ( .D(datain[5]), .E(n2359), .CK(clk), .QN(n2200) );
  EDFFX1 \img_buff_reg[58][4]  ( .D(datain[4]), .E(n2359), .CK(clk), .QN(n2166) );
  EDFFX1 \img_buff_reg[59][7]  ( .D(datain[7]), .E(n2358), .CK(clk), .QN(n2269) );
  EDFFX1 \img_buff_reg[59][6]  ( .D(datain[6]), .E(n2358), .CK(clk), .QN(n2235) );
  EDFFX1 \img_buff_reg[59][5]  ( .D(datain[5]), .E(n2358), .CK(clk), .QN(n2201) );
  EDFFX1 \img_buff_reg[59][4]  ( .D(datain[4]), .E(n2358), .CK(clk), .QN(n2167) );
  EDFFX1 \img_buff_reg[59][3]  ( .D(datain[3]), .E(n2358), .CK(clk), .QN(n2133) );
  EDFFX1 \img_buff_reg[59][2]  ( .D(datain[2]), .E(n2358), .CK(clk), .QN(n2099) );
  EDFFX1 \img_buff_reg[59][1]  ( .D(datain[1]), .E(n2358), .CK(clk), .QN(n2065) );
  EDFFX1 \img_buff_reg[59][0]  ( .D(datain[0]), .E(n2358), .CK(clk), .QN(n2031) );
  EDFFX1 \img_buff_reg[65][7]  ( .D(datain[7]), .E(n2352), .CK(clk), .QN(n328)
         );
  EDFFX1 \img_buff_reg[65][6]  ( .D(datain[6]), .E(n2352), .CK(clk), .QN(n329)
         );
  EDFFX1 \img_buff_reg[65][5]  ( .D(datain[5]), .E(n2352), .CK(clk), .QN(n330)
         );
  EDFFX1 \img_buff_reg[65][4]  ( .D(datain[4]), .E(n2352), .CK(clk), .QN(n331)
         );
  EDFFX1 \img_buff_reg[65][3]  ( .D(datain[3]), .E(n2352), .CK(clk), .QN(n332)
         );
  EDFFX1 \img_buff_reg[65][2]  ( .D(datain[2]), .E(n2352), .CK(clk), .QN(n333)
         );
  EDFFX1 \img_buff_reg[65][1]  ( .D(datain[1]), .E(n2352), .CK(clk), .QN(n334)
         );
  EDFFX1 \img_buff_reg[65][0]  ( .D(datain[0]), .E(n2352), .CK(clk), .QN(n335)
         );
  EDFFX1 \img_buff_reg[66][7]  ( .D(datain[7]), .E(n2351), .CK(clk), .QN(n336)
         );
  EDFFX1 \img_buff_reg[66][6]  ( .D(datain[6]), .E(n2351), .CK(clk), .QN(n337)
         );
  EDFFX1 \img_buff_reg[66][5]  ( .D(datain[5]), .E(n2351), .CK(clk), .QN(n338)
         );
  EDFFX1 \img_buff_reg[66][4]  ( .D(datain[4]), .E(n2351), .CK(clk), .QN(n339)
         );
  EDFFX1 \img_buff_reg[66][3]  ( .D(datain[3]), .E(n2351), .CK(clk), .QN(n340)
         );
  EDFFX1 \img_buff_reg[66][2]  ( .D(datain[2]), .E(n2351), .CK(clk), .QN(n341)
         );
  EDFFX1 \img_buff_reg[66][1]  ( .D(datain[1]), .E(n2351), .CK(clk), .QN(n342)
         );
  EDFFX1 \img_buff_reg[66][0]  ( .D(datain[0]), .E(n2351), .CK(clk), .QN(n343)
         );
  EDFFX1 \img_buff_reg[75][7]  ( .D(datain[7]), .E(n2342), .CK(clk), .QN(n2273) );
  EDFFX1 \img_buff_reg[75][6]  ( .D(datain[6]), .E(n2342), .CK(clk), .QN(n2239) );
  EDFFX1 \img_buff_reg[75][5]  ( .D(datain[5]), .E(n2342), .CK(clk), .QN(n2205) );
  EDFFX1 \img_buff_reg[75][4]  ( .D(datain[4]), .E(n2342), .CK(clk), .QN(n2171) );
  EDFFX1 \img_buff_reg[75][3]  ( .D(datain[3]), .E(n2342), .CK(clk), .QN(n2137) );
  EDFFX1 \img_buff_reg[75][2]  ( .D(datain[2]), .E(n2342), .CK(clk), .QN(n2103) );
  EDFFX1 \img_buff_reg[75][1]  ( .D(datain[1]), .E(n2342), .CK(clk), .QN(n2069) );
  EDFFX1 \img_buff_reg[75][0]  ( .D(datain[0]), .E(n2342), .CK(clk), .QN(n2035) );
  EDFFX1 \img_buff_reg[80][7]  ( .D(datain[7]), .E(n2337), .CK(clk), .QN(n2270) );
  EDFFX1 \img_buff_reg[80][6]  ( .D(datain[6]), .E(n2337), .CK(clk), .QN(n2236) );
  EDFFX1 \img_buff_reg[80][5]  ( .D(datain[5]), .E(n2337), .CK(clk), .QN(n2202) );
  EDFFX1 \img_buff_reg[80][4]  ( .D(datain[4]), .E(n2337), .CK(clk), .QN(n2168) );
  EDFFX1 \img_buff_reg[80][3]  ( .D(datain[3]), .E(n2337), .CK(clk), .QN(n2134) );
  EDFFX1 \img_buff_reg[80][2]  ( .D(datain[2]), .E(n2337), .CK(clk), .QN(n2100) );
  EDFFX1 \img_buff_reg[80][1]  ( .D(datain[1]), .E(n2337), .CK(clk), .QN(n2066) );
  EDFFX1 \img_buff_reg[80][0]  ( .D(datain[0]), .E(n2337), .CK(clk), .QN(n2032) );
  EDFFX1 \img_buff_reg[85][7]  ( .D(datain[7]), .E(n2332), .CK(clk), .QN(n2280) );
  EDFFX1 \img_buff_reg[85][6]  ( .D(datain[6]), .E(n2332), .CK(clk), .QN(n2246) );
  EDFFX1 \img_buff_reg[85][5]  ( .D(datain[5]), .E(n2332), .CK(clk), .QN(n2212) );
  EDFFX1 \img_buff_reg[85][4]  ( .D(datain[4]), .E(n2332), .CK(clk), .QN(n2178) );
  EDFFX1 \img_buff_reg[85][3]  ( .D(datain[3]), .E(n2332), .CK(clk), .QN(n2144) );
  EDFFX1 \img_buff_reg[85][2]  ( .D(datain[2]), .E(n2332), .CK(clk), .QN(n2110) );
  EDFFX1 \img_buff_reg[85][1]  ( .D(datain[1]), .E(n2332), .CK(clk), .QN(n2076) );
  EDFFX1 \img_buff_reg[85][0]  ( .D(datain[0]), .E(n2332), .CK(clk), .QN(n2042) );
  EDFFX1 \img_buff_reg[86][7]  ( .D(datain[7]), .E(n2331), .CK(clk), .QN(n2281) );
  EDFFX1 \img_buff_reg[86][6]  ( .D(datain[6]), .E(n2331), .CK(clk), .QN(n2247) );
  EDFFX1 \img_buff_reg[86][5]  ( .D(datain[5]), .E(n2331), .CK(clk), .QN(n2213) );
  EDFFX1 \img_buff_reg[86][4]  ( .D(datain[4]), .E(n2331), .CK(clk), .QN(n2179) );
  EDFFX1 \img_buff_reg[86][3]  ( .D(datain[3]), .E(n2331), .CK(clk), .QN(n2145) );
  EDFFX1 \img_buff_reg[86][2]  ( .D(datain[2]), .E(n2331), .CK(clk), .QN(n2111) );
  EDFFX1 \img_buff_reg[86][1]  ( .D(datain[1]), .E(n2331), .CK(clk), .QN(n2077) );
  EDFFX1 \img_buff_reg[86][0]  ( .D(datain[0]), .E(n2331), .CK(clk), .QN(n2043) );
  EDFFX1 \img_buff_reg[92][7]  ( .D(datain[7]), .E(n2325), .CK(clk), .QN(n2276) );
  EDFFX1 \img_buff_reg[92][6]  ( .D(datain[6]), .E(n2325), .CK(clk), .QN(n2242) );
  EDFFX1 \img_buff_reg[92][5]  ( .D(datain[5]), .E(n2325), .CK(clk), .QN(n2208) );
  EDFFX1 \img_buff_reg[92][4]  ( .D(datain[4]), .E(n2325), .CK(clk), .QN(n2174) );
  EDFFX1 \img_buff_reg[92][3]  ( .D(datain[3]), .E(n2325), .CK(clk), .QN(n2140) );
  EDFFX1 \img_buff_reg[92][2]  ( .D(datain[2]), .E(n2325), .CK(clk), .QN(n2106) );
  EDFFX1 \img_buff_reg[92][1]  ( .D(datain[1]), .E(n2325), .CK(clk), .QN(n2072) );
  EDFFX1 \img_buff_reg[92][0]  ( .D(datain[0]), .E(n2325), .CK(clk), .QN(n2038) );
  EDFFX1 \img_buff_reg[93][7]  ( .D(datain[7]), .E(n2324), .CK(clk), .QN(n2277) );
  EDFFX1 \img_buff_reg[93][6]  ( .D(datain[6]), .E(n2324), .CK(clk), .QN(n2243) );
  EDFFX1 \img_buff_reg[93][5]  ( .D(datain[5]), .E(n2324), .CK(clk), .QN(n2209) );
  EDFFX1 \img_buff_reg[93][4]  ( .D(datain[4]), .E(n2324), .CK(clk), .QN(n2175) );
  EDFFX1 \img_buff_reg[93][3]  ( .D(datain[3]), .E(n2324), .CK(clk), .QN(n2141) );
  EDFFX1 \img_buff_reg[93][2]  ( .D(datain[2]), .E(n2324), .CK(clk), .QN(n2107) );
  EDFFX1 \img_buff_reg[93][1]  ( .D(datain[1]), .E(n2324), .CK(clk), .QN(n2073) );
  EDFFX1 \img_buff_reg[93][0]  ( .D(datain[0]), .E(n2324), .CK(clk), .QN(n2039) );
  EDFFX1 \img_buff_reg[104][7]  ( .D(datain[7]), .E(n2313), .CK(clk), .QN(n408) );
  EDFFX1 \img_buff_reg[104][6]  ( .D(datain[6]), .E(n2313), .CK(clk), .QN(n409) );
  EDFFX1 \img_buff_reg[104][5]  ( .D(datain[5]), .E(n2313), .CK(clk), .QN(n410) );
  EDFFX1 \img_buff_reg[104][4]  ( .D(datain[4]), .E(n2313), .CK(clk), .QN(n411) );
  EDFFX1 \img_buff_reg[104][3]  ( .D(datain[3]), .E(n2313), .CK(clk), .QN(n412) );
  EDFFX1 \img_buff_reg[104][2]  ( .D(datain[2]), .E(n2313), .CK(clk), .QN(n413) );
  EDFFX1 \img_buff_reg[104][1]  ( .D(datain[1]), .E(n2313), .CK(clk), .QN(n414) );
  EDFFX1 \img_buff_reg[104][0]  ( .D(datain[0]), .E(n2313), .CK(clk), .QN(n415) );
  EDFFX1 \img_buff_reg[106][7]  ( .D(datain[7]), .E(n2311), .CK(clk), .QN(
        n2282) );
  EDFFX1 \img_buff_reg[106][6]  ( .D(datain[6]), .E(n2311), .CK(clk), .QN(
        n2248) );
  EDFFX1 \img_buff_reg[106][5]  ( .D(datain[5]), .E(n2311), .CK(clk), .QN(
        n2214) );
  EDFFX1 \img_buff_reg[106][4]  ( .D(datain[4]), .E(n2311), .CK(clk), .QN(
        n2180) );
  EDFFX1 \img_buff_reg[106][3]  ( .D(datain[3]), .E(n2311), .CK(clk), .QN(
        n2146) );
  EDFFX1 \img_buff_reg[106][2]  ( .D(datain[2]), .E(n2311), .CK(clk), .QN(
        n2112) );
  EDFFX1 \img_buff_reg[106][1]  ( .D(datain[1]), .E(n2311), .CK(clk), .QN(
        n2078) );
  EDFFX1 \img_buff_reg[106][0]  ( .D(datain[0]), .E(n2311), .CK(clk), .QN(
        n2044) );
  EDFFX1 \img_buff_reg[32][7]  ( .D(datain[7]), .E(n2385), .CK(clk), .QN(n2295) );
  EDFFX1 \img_buff_reg[32][6]  ( .D(datain[6]), .E(n2385), .CK(clk), .QN(n2261) );
  EDFFX1 \img_buff_reg[32][5]  ( .D(datain[5]), .E(n2385), .CK(clk), .QN(n2227) );
  EDFFX1 \img_buff_reg[32][4]  ( .D(datain[4]), .E(n2385), .CK(clk), .QN(n2193) );
  EDFFX1 \img_buff_reg[32][3]  ( .D(datain[3]), .E(n2385), .CK(clk), .QN(n2159) );
  EDFFX1 \img_buff_reg[32][2]  ( .D(datain[2]), .E(n2385), .CK(clk), .QN(n2125) );
  EDFFX1 \img_buff_reg[32][1]  ( .D(datain[1]), .E(n2385), .CK(clk), .QN(n2091) );
  EDFFX1 \img_buff_reg[32][0]  ( .D(datain[0]), .E(n2385), .CK(clk), .QN(n2057) );
  EDFFX1 \img_buff_reg[36][7]  ( .D(datain[7]), .E(n2381), .CK(clk), .QN(n280)
         );
  EDFFX1 \img_buff_reg[36][6]  ( .D(datain[6]), .E(n2381), .CK(clk), .QN(n281)
         );
  EDFFX1 \img_buff_reg[36][5]  ( .D(datain[5]), .E(n2381), .CK(clk), .QN(n282)
         );
  EDFFX1 \img_buff_reg[36][4]  ( .D(datain[4]), .E(n2381), .CK(clk), .QN(n283)
         );
  EDFFX1 \img_buff_reg[36][3]  ( .D(datain[3]), .E(n2381), .CK(clk), .QN(n284)
         );
  EDFFX1 \img_buff_reg[36][2]  ( .D(datain[2]), .E(n2381), .CK(clk), .QN(n285)
         );
  EDFFX1 \img_buff_reg[36][1]  ( .D(datain[1]), .E(n2381), .CK(clk), .QN(n286)
         );
  EDFFX1 \img_buff_reg[36][0]  ( .D(datain[0]), .E(n2381), .CK(clk), .QN(n287)
         );
  EDFFX1 \img_buff_reg[37][7]  ( .D(datain[7]), .E(n2380), .CK(clk), .QN(n288)
         );
  EDFFX1 \img_buff_reg[37][6]  ( .D(datain[6]), .E(n2380), .CK(clk), .QN(n289)
         );
  EDFFX1 \img_buff_reg[37][5]  ( .D(datain[5]), .E(n2380), .CK(clk), .QN(n290)
         );
  EDFFX1 \img_buff_reg[37][4]  ( .D(datain[4]), .E(n2380), .CK(clk), .QN(n291)
         );
  EDFFX1 \img_buff_reg[37][3]  ( .D(datain[3]), .E(n2380), .CK(clk), .QN(n292)
         );
  EDFFX1 \img_buff_reg[37][2]  ( .D(datain[2]), .E(n2380), .CK(clk), .QN(n293)
         );
  EDFFX1 \img_buff_reg[37][1]  ( .D(datain[1]), .E(n2380), .CK(clk), .QN(n294)
         );
  EDFFX1 \img_buff_reg[37][0]  ( .D(datain[0]), .E(n2380), .CK(clk), .QN(n295)
         );
  DFFSXL \W_reg[0]  ( .D(n1281), .CK(clk), .SN(n2309), .QN(n431) );
  DFFSXL \cmd_reg_reg[1]  ( .D(n1268), .CK(clk), .SN(n2309), .Q(n1282), .QN(
        n217) );
  DFFSXL \cmd_reg_reg[0]  ( .D(n1269), .CK(clk), .SN(n2309), .Q(n1285), .QN(
        n218) );
  DFFSXL \cmd_reg_reg[2]  ( .D(n1277), .CK(clk), .SN(n2309), .Q(n1283), .QN(
        n216) );
  DFFSXL \L_reg[1]  ( .D(n1264), .CK(clk), .SN(n2309), .QN(n426) );
  DFFSXL \L_reg[2]  ( .D(n1263), .CK(clk), .SN(n2309), .QN(n425) );
  DFFSXL \W_reg[2]  ( .D(n1279), .CK(clk), .SN(n2309), .QN(n429) );
  EDFFX1 \img_buff_reg[5][7]  ( .D(datain[7]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][7] ) );
  EDFFX1 \img_buff_reg[5][6]  ( .D(datain[6]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][6] ) );
  EDFFX1 \img_buff_reg[5][5]  ( .D(datain[5]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][5] ) );
  EDFFX1 \img_buff_reg[5][4]  ( .D(datain[4]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][4] ) );
  EDFFX1 \img_buff_reg[5][3]  ( .D(datain[3]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][3] ) );
  EDFFX1 \img_buff_reg[5][2]  ( .D(datain[2]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][2] ) );
  EDFFX1 \img_buff_reg[5][1]  ( .D(datain[1]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][1] ) );
  EDFFX1 \img_buff_reg[5][0]  ( .D(datain[0]), .E(n2412), .CK(clk), .Q(
        \img_buff[5][0] ) );
  EDFFX1 \img_buff_reg[12][7]  ( .D(datain[7]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][7] ) );
  EDFFX1 \img_buff_reg[12][6]  ( .D(datain[6]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][6] ) );
  EDFFX1 \img_buff_reg[12][5]  ( .D(datain[5]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][5] ) );
  EDFFX1 \img_buff_reg[12][4]  ( .D(datain[4]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][4] ) );
  EDFFX1 \img_buff_reg[12][3]  ( .D(datain[3]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][3] ) );
  EDFFX1 \img_buff_reg[12][2]  ( .D(datain[2]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][2] ) );
  EDFFX1 \img_buff_reg[12][1]  ( .D(datain[1]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][1] ) );
  EDFFX1 \img_buff_reg[12][0]  ( .D(datain[0]), .E(n2405), .CK(clk), .Q(
        \img_buff[12][0] ) );
  EDFFX1 \img_buff_reg[23][7]  ( .D(datain[7]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][7] ) );
  EDFFX1 \img_buff_reg[23][6]  ( .D(datain[6]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][6] ) );
  EDFFX1 \img_buff_reg[23][5]  ( .D(datain[5]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][5] ) );
  EDFFX1 \img_buff_reg[23][4]  ( .D(datain[4]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][4] ) );
  EDFFX1 \img_buff_reg[23][3]  ( .D(datain[3]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][3] ) );
  EDFFX1 \img_buff_reg[23][2]  ( .D(datain[2]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][2] ) );
  EDFFX1 \img_buff_reg[23][1]  ( .D(datain[1]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][1] ) );
  EDFFX1 \img_buff_reg[23][0]  ( .D(datain[0]), .E(n2394), .CK(clk), .Q(
        \img_buff[23][0] ) );
  EDFFX1 \img_buff_reg[28][7]  ( .D(datain[7]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][7] ) );
  EDFFX1 \img_buff_reg[28][6]  ( .D(datain[6]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][6] ) );
  EDFFX1 \img_buff_reg[28][5]  ( .D(datain[5]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][5] ) );
  EDFFX1 \img_buff_reg[28][4]  ( .D(datain[4]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][4] ) );
  EDFFX1 \img_buff_reg[28][3]  ( .D(datain[3]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][3] ) );
  EDFFX1 \img_buff_reg[28][2]  ( .D(datain[2]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][2] ) );
  EDFFX1 \img_buff_reg[28][1]  ( .D(datain[1]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][1] ) );
  EDFFX1 \img_buff_reg[28][0]  ( .D(datain[0]), .E(n2389), .CK(clk), .Q(
        \img_buff[28][0] ) );
  EDFFX1 \img_buff_reg[50][7]  ( .D(datain[7]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][7] ) );
  EDFFX1 \img_buff_reg[50][6]  ( .D(datain[6]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][6] ) );
  EDFFX1 \img_buff_reg[50][5]  ( .D(datain[5]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][5] ) );
  EDFFX1 \img_buff_reg[50][4]  ( .D(datain[4]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][4] ) );
  EDFFX1 \img_buff_reg[50][3]  ( .D(datain[3]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][3] ) );
  EDFFX1 \img_buff_reg[50][2]  ( .D(datain[2]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][2] ) );
  EDFFX1 \img_buff_reg[50][1]  ( .D(datain[1]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][1] ) );
  EDFFX1 \img_buff_reg[50][0]  ( .D(datain[0]), .E(n2367), .CK(clk), .Q(
        \img_buff[50][0] ) );
  EDFFX1 \img_buff_reg[55][7]  ( .D(datain[7]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][7] ) );
  EDFFX1 \img_buff_reg[55][6]  ( .D(datain[6]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][6] ) );
  EDFFX1 \img_buff_reg[55][5]  ( .D(datain[5]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][5] ) );
  EDFFX1 \img_buff_reg[55][4]  ( .D(datain[4]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][4] ) );
  EDFFX1 \img_buff_reg[55][3]  ( .D(datain[3]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][3] ) );
  EDFFX1 \img_buff_reg[55][2]  ( .D(datain[2]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][2] ) );
  EDFFX1 \img_buff_reg[55][1]  ( .D(datain[1]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][1] ) );
  EDFFX1 \img_buff_reg[55][0]  ( .D(datain[0]), .E(n2362), .CK(clk), .Q(
        \img_buff[55][0] ) );
  EDFFX1 \img_buff_reg[64][7]  ( .D(datain[7]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][7] ) );
  EDFFX1 \img_buff_reg[64][6]  ( .D(datain[6]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][6] ) );
  EDFFX1 \img_buff_reg[64][5]  ( .D(datain[5]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][5] ) );
  EDFFX1 \img_buff_reg[64][4]  ( .D(datain[4]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][4] ) );
  EDFFX1 \img_buff_reg[64][3]  ( .D(datain[3]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][3] ) );
  EDFFX1 \img_buff_reg[64][2]  ( .D(datain[2]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][2] ) );
  EDFFX1 \img_buff_reg[64][1]  ( .D(datain[1]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][1] ) );
  EDFFX1 \img_buff_reg[64][0]  ( .D(datain[0]), .E(n2353), .CK(clk), .Q(
        \img_buff[64][0] ) );
  EDFFX1 \img_buff_reg[79][7]  ( .D(datain[7]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][7] ) );
  EDFFX1 \img_buff_reg[79][6]  ( .D(datain[6]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][6] ) );
  EDFFX1 \img_buff_reg[79][5]  ( .D(datain[5]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][5] ) );
  EDFFX1 \img_buff_reg[79][4]  ( .D(datain[4]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][4] ) );
  EDFFX1 \img_buff_reg[79][3]  ( .D(datain[3]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][3] ) );
  EDFFX1 \img_buff_reg[79][2]  ( .D(datain[2]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][2] ) );
  EDFFX1 \img_buff_reg[79][1]  ( .D(datain[1]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][1] ) );
  EDFFX1 \img_buff_reg[79][0]  ( .D(datain[0]), .E(n2338), .CK(clk), .Q(
        \img_buff[79][0] ) );
  EDFFX1 \img_buff_reg[82][7]  ( .D(datain[7]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][7] ) );
  EDFFX1 \img_buff_reg[82][6]  ( .D(datain[6]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][6] ) );
  EDFFX1 \img_buff_reg[82][5]  ( .D(datain[5]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][5] ) );
  EDFFX1 \img_buff_reg[82][4]  ( .D(datain[4]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][4] ) );
  EDFFX1 \img_buff_reg[82][3]  ( .D(datain[3]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][3] ) );
  EDFFX1 \img_buff_reg[82][2]  ( .D(datain[2]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][2] ) );
  EDFFX1 \img_buff_reg[82][1]  ( .D(datain[1]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][1] ) );
  EDFFX1 \img_buff_reg[82][0]  ( .D(datain[0]), .E(n2335), .CK(clk), .Q(
        \img_buff[82][0] ) );
  EDFFX1 \img_buff_reg[102][7]  ( .D(datain[7]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][7] ) );
  EDFFX1 \img_buff_reg[102][6]  ( .D(datain[6]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][6] ) );
  EDFFX1 \img_buff_reg[102][5]  ( .D(datain[5]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][5] ) );
  EDFFX1 \img_buff_reg[102][4]  ( .D(datain[4]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][4] ) );
  EDFFX1 \img_buff_reg[102][3]  ( .D(datain[3]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][3] ) );
  EDFFX1 \img_buff_reg[102][2]  ( .D(datain[2]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][2] ) );
  EDFFX1 \img_buff_reg[102][1]  ( .D(datain[1]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][1] ) );
  EDFFX1 \img_buff_reg[102][0]  ( .D(datain[0]), .E(n2315), .CK(clk), .Q(
        \img_buff[102][0] ) );
  EDFFX1 \img_buff_reg[39][7]  ( .D(datain[7]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][7] ) );
  EDFFX1 \img_buff_reg[39][6]  ( .D(datain[6]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][6] ) );
  EDFFX1 \img_buff_reg[39][5]  ( .D(datain[5]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][5] ) );
  EDFFX1 \img_buff_reg[39][4]  ( .D(datain[4]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][4] ) );
  EDFFX1 \img_buff_reg[39][3]  ( .D(datain[3]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][3] ) );
  EDFFX1 \img_buff_reg[39][2]  ( .D(datain[2]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][2] ) );
  EDFFX1 \img_buff_reg[39][1]  ( .D(datain[1]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][1] ) );
  EDFFX1 \img_buff_reg[39][0]  ( .D(datain[0]), .E(n2378), .CK(clk), .Q(
        \img_buff[39][0] ) );
  EDFFX1 \img_buff_reg[19][7]  ( .D(datain[7]), .E(n2398), .CK(clk), .Q(n2292)
         );
  EDFFX1 \img_buff_reg[19][6]  ( .D(datain[6]), .E(n2398), .CK(clk), .Q(n2258)
         );
  EDFFX1 \img_buff_reg[19][5]  ( .D(datain[5]), .E(n2398), .CK(clk), .Q(n2224)
         );
  EDFFX1 \img_buff_reg[19][4]  ( .D(datain[4]), .E(n2398), .CK(clk), .Q(n2190)
         );
  EDFFX1 \img_buff_reg[19][3]  ( .D(datain[3]), .E(n2398), .CK(clk), .Q(n2156)
         );
  EDFFX1 \img_buff_reg[19][2]  ( .D(datain[2]), .E(n2398), .CK(clk), .Q(n2122)
         );
  EDFFX1 \img_buff_reg[19][1]  ( .D(datain[1]), .E(n2398), .CK(clk), .Q(n2088)
         );
  EDFFX1 \img_buff_reg[19][0]  ( .D(datain[0]), .E(n2398), .CK(clk), .Q(n2054)
         );
  EDFFX1 \img_buff_reg[25][7]  ( .D(datain[7]), .E(n2392), .CK(clk), .Q(n2290)
         );
  EDFFX1 \img_buff_reg[25][6]  ( .D(datain[6]), .E(n2392), .CK(clk), .Q(n2256)
         );
  EDFFX1 \img_buff_reg[25][5]  ( .D(datain[5]), .E(n2392), .CK(clk), .Q(n2222)
         );
  EDFFX1 \img_buff_reg[25][4]  ( .D(datain[4]), .E(n2392), .CK(clk), .Q(n2188)
         );
  EDFFX1 \img_buff_reg[25][3]  ( .D(datain[3]), .E(n2392), .CK(clk), .Q(n2154)
         );
  EDFFX1 \img_buff_reg[25][2]  ( .D(datain[2]), .E(n2392), .CK(clk), .Q(n2120)
         );
  EDFFX1 \img_buff_reg[25][1]  ( .D(datain[1]), .E(n2392), .CK(clk), .Q(n2086)
         );
  EDFFX1 \img_buff_reg[25][0]  ( .D(datain[0]), .E(n2392), .CK(clk), .Q(n2052)
         );
  EDFFX1 \img_buff_reg[26][7]  ( .D(datain[7]), .E(n2391), .CK(clk), .Q(n2289)
         );
  EDFFX1 \img_buff_reg[26][6]  ( .D(datain[6]), .E(n2391), .CK(clk), .Q(n2255)
         );
  EDFFX1 \img_buff_reg[26][5]  ( .D(datain[5]), .E(n2391), .CK(clk), .Q(n2221)
         );
  EDFFX1 \img_buff_reg[26][4]  ( .D(datain[4]), .E(n2391), .CK(clk), .Q(n2187)
         );
  EDFFX1 \img_buff_reg[26][3]  ( .D(datain[3]), .E(n2391), .CK(clk), .Q(n2153)
         );
  EDFFX1 \img_buff_reg[26][2]  ( .D(datain[2]), .E(n2391), .CK(clk), .Q(n2119)
         );
  EDFFX1 \img_buff_reg[26][1]  ( .D(datain[1]), .E(n2391), .CK(clk), .Q(n2085)
         );
  EDFFX1 \img_buff_reg[26][0]  ( .D(datain[0]), .E(n2391), .CK(clk), .Q(n2051)
         );
  EDFFX1 \img_buff_reg[52][7]  ( .D(datain[7]), .E(n2365), .CK(clk), .Q(n2298)
         );
  EDFFX1 \img_buff_reg[52][6]  ( .D(datain[6]), .E(n2365), .CK(clk), .Q(n2264)
         );
  EDFFX1 \img_buff_reg[52][5]  ( .D(datain[5]), .E(n2365), .CK(clk), .Q(n2230)
         );
  EDFFX1 \img_buff_reg[52][4]  ( .D(datain[4]), .E(n2365), .CK(clk), .Q(n2196)
         );
  EDFFX1 \img_buff_reg[52][3]  ( .D(datain[3]), .E(n2365), .CK(clk), .Q(n2162)
         );
  EDFFX1 \img_buff_reg[52][2]  ( .D(datain[2]), .E(n2365), .CK(clk), .Q(n2128)
         );
  EDFFX1 \img_buff_reg[52][1]  ( .D(datain[1]), .E(n2365), .CK(clk), .Q(n2094)
         );
  EDFFX1 \img_buff_reg[52][0]  ( .D(datain[0]), .E(n2365), .CK(clk), .Q(n2060)
         );
  EDFFX1 \img_buff_reg[53][7]  ( .D(datain[7]), .E(n2364), .CK(clk), .Q(n2297)
         );
  EDFFX1 \img_buff_reg[53][6]  ( .D(datain[6]), .E(n2364), .CK(clk), .Q(n2263)
         );
  EDFFX1 \img_buff_reg[53][5]  ( .D(datain[5]), .E(n2364), .CK(clk), .Q(n2229)
         );
  EDFFX1 \img_buff_reg[53][4]  ( .D(datain[4]), .E(n2364), .CK(clk), .Q(n2195)
         );
  EDFFX1 \img_buff_reg[53][3]  ( .D(datain[3]), .E(n2364), .CK(clk), .Q(n2161)
         );
  EDFFX1 \img_buff_reg[53][2]  ( .D(datain[2]), .E(n2364), .CK(clk), .Q(n2127)
         );
  EDFFX1 \img_buff_reg[53][1]  ( .D(datain[1]), .E(n2364), .CK(clk), .Q(n2093)
         );
  EDFFX1 \img_buff_reg[53][0]  ( .D(datain[0]), .E(n2364), .CK(clk), .Q(n2059)
         );
  EDFFX1 \img_buff_reg[71][7]  ( .D(datain[7]), .E(n2346), .CK(clk), .Q(n2274)
         );
  EDFFX1 \img_buff_reg[71][6]  ( .D(datain[6]), .E(n2346), .CK(clk), .Q(n2240)
         );
  EDFFX1 \img_buff_reg[71][5]  ( .D(datain[5]), .E(n2346), .CK(clk), .Q(n2206)
         );
  EDFFX1 \img_buff_reg[71][4]  ( .D(datain[4]), .E(n2346), .CK(clk), .Q(n2172)
         );
  EDFFX1 \img_buff_reg[71][3]  ( .D(datain[3]), .E(n2346), .CK(clk), .Q(n2138)
         );
  EDFFX1 \img_buff_reg[71][2]  ( .D(datain[2]), .E(n2346), .CK(clk), .Q(n2104)
         );
  EDFFX1 \img_buff_reg[71][1]  ( .D(datain[1]), .E(n2346), .CK(clk), .Q(n2070)
         );
  EDFFX1 \img_buff_reg[71][0]  ( .D(datain[0]), .E(n2346), .CK(clk), .Q(n2036)
         );
  EDFFX1 \img_buff_reg[77][7]  ( .D(datain[7]), .E(n2340), .CK(clk), .Q(n2272)
         );
  EDFFX1 \img_buff_reg[77][6]  ( .D(datain[6]), .E(n2340), .CK(clk), .Q(n2238)
         );
  EDFFX1 \img_buff_reg[77][5]  ( .D(datain[5]), .E(n2340), .CK(clk), .Q(n2204)
         );
  EDFFX1 \img_buff_reg[77][4]  ( .D(datain[4]), .E(n2340), .CK(clk), .Q(n2170)
         );
  EDFFX1 \img_buff_reg[77][3]  ( .D(datain[3]), .E(n2340), .CK(clk), .Q(n2136)
         );
  EDFFX1 \img_buff_reg[77][2]  ( .D(datain[2]), .E(n2340), .CK(clk), .Q(n2102)
         );
  EDFFX1 \img_buff_reg[77][1]  ( .D(datain[1]), .E(n2340), .CK(clk), .Q(n2068)
         );
  EDFFX1 \img_buff_reg[77][0]  ( .D(datain[0]), .E(n2340), .CK(clk), .Q(n2034)
         );
  EDFFX1 \img_buff_reg[78][7]  ( .D(datain[7]), .E(n2339), .CK(clk), .Q(n2271)
         );
  EDFFX1 \img_buff_reg[78][6]  ( .D(datain[6]), .E(n2339), .CK(clk), .Q(n2237)
         );
  EDFFX1 \img_buff_reg[78][5]  ( .D(datain[5]), .E(n2339), .CK(clk), .Q(n2203)
         );
  EDFFX1 \img_buff_reg[78][4]  ( .D(datain[4]), .E(n2339), .CK(clk), .Q(n2169)
         );
  EDFFX1 \img_buff_reg[78][3]  ( .D(datain[3]), .E(n2339), .CK(clk), .Q(n2135)
         );
  EDFFX1 \img_buff_reg[78][2]  ( .D(datain[2]), .E(n2339), .CK(clk), .Q(n2101)
         );
  EDFFX1 \img_buff_reg[78][1]  ( .D(datain[1]), .E(n2339), .CK(clk), .Q(n2067)
         );
  EDFFX1 \img_buff_reg[78][0]  ( .D(datain[0]), .E(n2339), .CK(clk), .Q(n2033)
         );
  EDFFX1 \img_buff_reg[91][7]  ( .D(datain[7]), .E(n2326), .CK(clk), .Q(n2278)
         );
  EDFFX1 \img_buff_reg[91][6]  ( .D(datain[6]), .E(n2326), .CK(clk), .Q(n2244)
         );
  EDFFX1 \img_buff_reg[91][5]  ( .D(datain[5]), .E(n2326), .CK(clk), .Q(n2210)
         );
  EDFFX1 \img_buff_reg[91][4]  ( .D(datain[4]), .E(n2326), .CK(clk), .Q(n2176)
         );
  EDFFX1 \img_buff_reg[91][3]  ( .D(datain[3]), .E(n2326), .CK(clk), .Q(n2142)
         );
  EDFFX1 \img_buff_reg[91][2]  ( .D(datain[2]), .E(n2326), .CK(clk), .Q(n2108)
         );
  EDFFX1 \img_buff_reg[91][1]  ( .D(datain[1]), .E(n2326), .CK(clk), .Q(n2074)
         );
  EDFFX1 \img_buff_reg[91][0]  ( .D(datain[0]), .E(n2326), .CK(clk), .Q(n2040)
         );
  EDFFX1 \img_buff_reg[100][7]  ( .D(datain[7]), .E(n2317), .CK(clk), .Q(n2284) );
  EDFFX1 \img_buff_reg[100][6]  ( .D(datain[6]), .E(n2317), .CK(clk), .Q(n2250) );
  EDFFX1 \img_buff_reg[100][5]  ( .D(datain[5]), .E(n2317), .CK(clk), .Q(n2216) );
  EDFFX1 \img_buff_reg[100][4]  ( .D(datain[4]), .E(n2317), .CK(clk), .Q(n2182) );
  EDFFX1 \img_buff_reg[100][3]  ( .D(datain[3]), .E(n2317), .CK(clk), .Q(n2148) );
  EDFFX1 \img_buff_reg[100][2]  ( .D(datain[2]), .E(n2317), .CK(clk), .Q(n2114) );
  EDFFX1 \img_buff_reg[100][1]  ( .D(datain[1]), .E(n2317), .CK(clk), .Q(n2080) );
  EDFFX1 \img_buff_reg[100][0]  ( .D(datain[0]), .E(n2317), .CK(clk), .Q(n2046) );
  EDFFX1 \img_buff_reg[105][7]  ( .D(datain[7]), .E(n2312), .CK(clk), .Q(n2283) );
  EDFFX1 \img_buff_reg[105][6]  ( .D(datain[6]), .E(n2312), .CK(clk), .Q(n2249) );
  EDFFX1 \img_buff_reg[105][5]  ( .D(datain[5]), .E(n2312), .CK(clk), .Q(n2215) );
  EDFFX1 \img_buff_reg[105][4]  ( .D(datain[4]), .E(n2312), .CK(clk), .Q(n2181) );
  EDFFX1 \img_buff_reg[105][3]  ( .D(datain[3]), .E(n2312), .CK(clk), .Q(n2147) );
  EDFFX1 \img_buff_reg[105][2]  ( .D(datain[2]), .E(n2312), .CK(clk), .Q(n2113) );
  EDFFX1 \img_buff_reg[105][1]  ( .D(datain[1]), .E(n2312), .CK(clk), .Q(n2079) );
  EDFFX1 \img_buff_reg[105][0]  ( .D(datain[0]), .E(n2312), .CK(clk), .Q(n2045) );
  EDFFX1 \img_buff_reg[46][6]  ( .D(datain[6]), .E(n2371), .CK(clk), .Q(n2266)
         );
  EDFFX1 \img_buff_reg[46][5]  ( .D(datain[5]), .E(n2371), .CK(clk), .Q(n2232)
         );
  EDFFX1 \img_buff_reg[46][4]  ( .D(datain[4]), .E(n2371), .CK(clk), .Q(n2198)
         );
  EDFFX1 \img_buff_reg[46][3]  ( .D(datain[3]), .E(n2371), .CK(clk), .Q(n2164)
         );
  EDFFX1 \img_buff_reg[46][2]  ( .D(datain[2]), .E(n2371), .CK(clk), .Q(n2130)
         );
  EDFFX1 \img_buff_reg[46][1]  ( .D(datain[1]), .E(n2371), .CK(clk), .Q(n2096)
         );
  EDFFX1 \img_buff_reg[46][0]  ( .D(datain[0]), .E(n2371), .CK(clk), .Q(n2062)
         );
  EDFFX1 \img_buff_reg[46][7]  ( .D(datain[7]), .E(n2371), .CK(clk), .Q(n2300)
         );
  EDFFX1 \img_buff_reg[4][7]  ( .D(datain[7]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][7] ) );
  EDFFX1 \img_buff_reg[4][6]  ( .D(datain[6]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][6] ) );
  EDFFX1 \img_buff_reg[4][5]  ( .D(datain[5]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][5] ) );
  EDFFX1 \img_buff_reg[4][4]  ( .D(datain[4]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][4] ) );
  EDFFX1 \img_buff_reg[4][3]  ( .D(datain[3]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][3] ) );
  EDFFX1 \img_buff_reg[4][2]  ( .D(datain[2]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][2] ) );
  EDFFX1 \img_buff_reg[4][1]  ( .D(datain[1]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][1] ) );
  EDFFX1 \img_buff_reg[4][0]  ( .D(datain[0]), .E(n2413), .CK(clk), .Q(
        \img_buff[4][0] ) );
  EDFFX1 \img_buff_reg[11][7]  ( .D(datain[7]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][7] ) );
  EDFFX1 \img_buff_reg[11][6]  ( .D(datain[6]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][6] ) );
  EDFFX1 \img_buff_reg[11][5]  ( .D(datain[5]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][5] ) );
  EDFFX1 \img_buff_reg[11][4]  ( .D(datain[4]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][4] ) );
  EDFFX1 \img_buff_reg[11][3]  ( .D(datain[3]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][3] ) );
  EDFFX1 \img_buff_reg[11][2]  ( .D(datain[2]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][2] ) );
  EDFFX1 \img_buff_reg[11][1]  ( .D(datain[1]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][1] ) );
  EDFFX1 \img_buff_reg[11][0]  ( .D(datain[0]), .E(n2406), .CK(clk), .Q(
        \img_buff[11][0] ) );
  EDFFX1 \img_buff_reg[30][7]  ( .D(datain[7]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][7] ) );
  EDFFX1 \img_buff_reg[30][6]  ( .D(datain[6]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][6] ) );
  EDFFX1 \img_buff_reg[30][5]  ( .D(datain[5]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][5] ) );
  EDFFX1 \img_buff_reg[30][4]  ( .D(datain[4]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][4] ) );
  EDFFX1 \img_buff_reg[30][3]  ( .D(datain[3]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][3] ) );
  EDFFX1 \img_buff_reg[30][2]  ( .D(datain[2]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][2] ) );
  EDFFX1 \img_buff_reg[30][1]  ( .D(datain[1]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][1] ) );
  EDFFX1 \img_buff_reg[30][0]  ( .D(datain[0]), .E(n2387), .CK(clk), .Q(
        \img_buff[30][0] ) );
  EDFFX1 \img_buff_reg[57][7]  ( .D(datain[7]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][7] ) );
  EDFFX1 \img_buff_reg[57][6]  ( .D(datain[6]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][6] ) );
  EDFFX1 \img_buff_reg[57][5]  ( .D(datain[5]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][5] ) );
  EDFFX1 \img_buff_reg[57][4]  ( .D(datain[4]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][4] ) );
  EDFFX1 \img_buff_reg[57][3]  ( .D(datain[3]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][3] ) );
  EDFFX1 \img_buff_reg[57][2]  ( .D(datain[2]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][2] ) );
  EDFFX1 \img_buff_reg[57][1]  ( .D(datain[1]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][1] ) );
  EDFFX1 \img_buff_reg[57][0]  ( .D(datain[0]), .E(n2360), .CK(clk), .Q(
        \img_buff[57][0] ) );
  EDFFX1 \img_buff_reg[63][7]  ( .D(datain[7]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][7] ) );
  EDFFX1 \img_buff_reg[63][6]  ( .D(datain[6]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][6] ) );
  EDFFX1 \img_buff_reg[63][5]  ( .D(datain[5]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][5] ) );
  EDFFX1 \img_buff_reg[63][4]  ( .D(datain[4]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][4] ) );
  EDFFX1 \img_buff_reg[63][3]  ( .D(datain[3]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][3] ) );
  EDFFX1 \img_buff_reg[63][2]  ( .D(datain[2]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][2] ) );
  EDFFX1 \img_buff_reg[63][1]  ( .D(datain[1]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][1] ) );
  EDFFX1 \img_buff_reg[63][0]  ( .D(datain[0]), .E(n2354), .CK(clk), .Q(
        \img_buff[63][0] ) );
  EDFFX1 \img_buff_reg[84][7]  ( .D(datain[7]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][7] ) );
  EDFFX1 \img_buff_reg[84][6]  ( .D(datain[6]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][6] ) );
  EDFFX1 \img_buff_reg[84][5]  ( .D(datain[5]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][5] ) );
  EDFFX1 \img_buff_reg[84][4]  ( .D(datain[4]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][4] ) );
  EDFFX1 \img_buff_reg[84][3]  ( .D(datain[3]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][3] ) );
  EDFFX1 \img_buff_reg[84][2]  ( .D(datain[2]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][2] ) );
  EDFFX1 \img_buff_reg[84][1]  ( .D(datain[1]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][1] ) );
  EDFFX1 \img_buff_reg[84][0]  ( .D(datain[0]), .E(n2333), .CK(clk), .Q(
        \img_buff[84][0] ) );
  EDFFX1 \img_buff_reg[107][7]  ( .D(datain[7]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][7] ) );
  EDFFX1 \img_buff_reg[107][6]  ( .D(datain[6]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][6] ) );
  EDFFX1 \img_buff_reg[107][5]  ( .D(datain[5]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][5] ) );
  EDFFX1 \img_buff_reg[107][4]  ( .D(datain[4]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][4] ) );
  EDFFX1 \img_buff_reg[107][3]  ( .D(datain[3]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][3] ) );
  EDFFX1 \img_buff_reg[107][2]  ( .D(datain[2]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][2] ) );
  EDFFX1 \img_buff_reg[107][1]  ( .D(datain[1]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][1] ) );
  EDFFX1 \img_buff_reg[107][0]  ( .D(datain[0]), .E(n2310), .CK(clk), .Q(
        \img_buff[107][0] ) );
  EDFFX1 \img_buff_reg[38][7]  ( .D(datain[7]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][7] ) );
  EDFFX1 \img_buff_reg[38][6]  ( .D(datain[6]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][6] ) );
  EDFFX1 \img_buff_reg[38][5]  ( .D(datain[5]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][5] ) );
  EDFFX1 \img_buff_reg[38][4]  ( .D(datain[4]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][4] ) );
  EDFFX1 \img_buff_reg[38][3]  ( .D(datain[3]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][3] ) );
  EDFFX1 \img_buff_reg[38][2]  ( .D(datain[2]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][2] ) );
  EDFFX1 \img_buff_reg[38][1]  ( .D(datain[1]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][1] ) );
  EDFFX1 \img_buff_reg[38][0]  ( .D(datain[0]), .E(n2379), .CK(clk), .Q(
        \img_buff[38][0] ) );
  EDFFX1 \img_buff_reg[90][7]  ( .D(datain[7]), .E(n2327), .CK(clk), .Q(n2279)
         );
  EDFFX1 \img_buff_reg[90][6]  ( .D(datain[6]), .E(n2327), .CK(clk), .Q(n2245)
         );
  EDFFX1 \img_buff_reg[90][5]  ( .D(datain[5]), .E(n2327), .CK(clk), .Q(n2211)
         );
  EDFFX1 \img_buff_reg[90][4]  ( .D(datain[4]), .E(n2327), .CK(clk), .Q(n2177)
         );
  EDFFX1 \img_buff_reg[90][3]  ( .D(datain[3]), .E(n2327), .CK(clk), .Q(n2143)
         );
  EDFFX1 \img_buff_reg[90][2]  ( .D(datain[2]), .E(n2327), .CK(clk), .Q(n2109)
         );
  EDFFX1 \img_buff_reg[90][1]  ( .D(datain[1]), .E(n2327), .CK(clk), .Q(n2075)
         );
  EDFFX1 \img_buff_reg[90][0]  ( .D(datain[0]), .E(n2327), .CK(clk), .Q(n2041)
         );
  EDFFX1 \img_buff_reg[0][7]  ( .D(datain[7]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][7] ) );
  EDFFX1 \img_buff_reg[0][6]  ( .D(datain[6]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][6] ) );
  EDFFX1 \img_buff_reg[0][5]  ( .D(datain[5]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][5] ) );
  EDFFX1 \img_buff_reg[0][4]  ( .D(datain[4]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][4] ) );
  EDFFX1 \img_buff_reg[0][3]  ( .D(datain[3]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][3] ) );
  EDFFX1 \img_buff_reg[0][2]  ( .D(datain[2]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][2] ) );
  EDFFX1 \img_buff_reg[0][1]  ( .D(datain[1]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][1] ) );
  EDFFX1 \img_buff_reg[0][0]  ( .D(datain[0]), .E(n2417), .CK(clk), .Q(
        \img_buff[0][0] ) );
  EDFFX1 \img_buff_reg[8][7]  ( .D(datain[7]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][7] ) );
  EDFFX1 \img_buff_reg[8][6]  ( .D(datain[6]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][6] ) );
  EDFFX1 \img_buff_reg[8][5]  ( .D(datain[5]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][5] ) );
  EDFFX1 \img_buff_reg[8][4]  ( .D(datain[4]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][4] ) );
  EDFFX1 \img_buff_reg[8][3]  ( .D(datain[3]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][3] ) );
  EDFFX1 \img_buff_reg[8][2]  ( .D(datain[2]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][2] ) );
  EDFFX1 \img_buff_reg[8][1]  ( .D(datain[1]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][1] ) );
  EDFFX1 \img_buff_reg[8][0]  ( .D(datain[0]), .E(n2409), .CK(clk), .Q(
        \img_buff[8][0] ) );
  EDFFX1 \img_buff_reg[15][7]  ( .D(datain[7]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][7] ) );
  EDFFX1 \img_buff_reg[15][6]  ( .D(datain[6]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][6] ) );
  EDFFX1 \img_buff_reg[15][5]  ( .D(datain[5]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][5] ) );
  EDFFX1 \img_buff_reg[15][4]  ( .D(datain[4]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][4] ) );
  EDFFX1 \img_buff_reg[15][3]  ( .D(datain[3]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][3] ) );
  EDFFX1 \img_buff_reg[15][2]  ( .D(datain[2]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][2] ) );
  EDFFX1 \img_buff_reg[15][1]  ( .D(datain[1]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][1] ) );
  EDFFX1 \img_buff_reg[15][0]  ( .D(datain[0]), .E(n2402), .CK(clk), .Q(
        \img_buff[15][0] ) );
  EDFFX1 \img_buff_reg[16][7]  ( .D(datain[7]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][7] ) );
  EDFFX1 \img_buff_reg[16][6]  ( .D(datain[6]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][6] ) );
  EDFFX1 \img_buff_reg[16][5]  ( .D(datain[5]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][5] ) );
  EDFFX1 \img_buff_reg[16][4]  ( .D(datain[4]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][4] ) );
  EDFFX1 \img_buff_reg[16][3]  ( .D(datain[3]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][3] ) );
  EDFFX1 \img_buff_reg[16][2]  ( .D(datain[2]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][2] ) );
  EDFFX1 \img_buff_reg[16][1]  ( .D(datain[1]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][1] ) );
  EDFFX1 \img_buff_reg[16][0]  ( .D(datain[0]), .E(n2401), .CK(clk), .Q(
        \img_buff[16][0] ) );
  EDFFX1 \img_buff_reg[20][7]  ( .D(datain[7]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][7] ) );
  EDFFX1 \img_buff_reg[20][6]  ( .D(datain[6]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][6] ) );
  EDFFX1 \img_buff_reg[20][5]  ( .D(datain[5]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][5] ) );
  EDFFX1 \img_buff_reg[20][4]  ( .D(datain[4]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][4] ) );
  EDFFX1 \img_buff_reg[20][3]  ( .D(datain[3]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][3] ) );
  EDFFX1 \img_buff_reg[20][2]  ( .D(datain[2]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][2] ) );
  EDFFX1 \img_buff_reg[20][1]  ( .D(datain[1]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][1] ) );
  EDFFX1 \img_buff_reg[20][0]  ( .D(datain[0]), .E(n2397), .CK(clk), .Q(
        \img_buff[20][0] ) );
  EDFFX1 \img_buff_reg[27][7]  ( .D(datain[7]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][7] ) );
  EDFFX1 \img_buff_reg[27][6]  ( .D(datain[6]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][6] ) );
  EDFFX1 \img_buff_reg[27][5]  ( .D(datain[5]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][5] ) );
  EDFFX1 \img_buff_reg[27][4]  ( .D(datain[4]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][4] ) );
  EDFFX1 \img_buff_reg[27][3]  ( .D(datain[3]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][3] ) );
  EDFFX1 \img_buff_reg[27][2]  ( .D(datain[2]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][2] ) );
  EDFFX1 \img_buff_reg[27][1]  ( .D(datain[1]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][1] ) );
  EDFFX1 \img_buff_reg[27][0]  ( .D(datain[0]), .E(n2390), .CK(clk), .Q(
        \img_buff[27][0] ) );
  EDFFX1 \img_buff_reg[54][7]  ( .D(datain[7]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][7] ) );
  EDFFX1 \img_buff_reg[54][6]  ( .D(datain[6]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][6] ) );
  EDFFX1 \img_buff_reg[54][5]  ( .D(datain[5]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][5] ) );
  EDFFX1 \img_buff_reg[54][4]  ( .D(datain[4]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][4] ) );
  EDFFX1 \img_buff_reg[54][3]  ( .D(datain[3]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][3] ) );
  EDFFX1 \img_buff_reg[54][2]  ( .D(datain[2]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][2] ) );
  EDFFX1 \img_buff_reg[54][1]  ( .D(datain[1]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][1] ) );
  EDFFX1 \img_buff_reg[54][0]  ( .D(datain[0]), .E(n2363), .CK(clk), .Q(
        \img_buff[54][0] ) );
  EDFFX1 \img_buff_reg[62][7]  ( .D(datain[7]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][7] ) );
  EDFFX1 \img_buff_reg[62][6]  ( .D(datain[6]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][6] ) );
  EDFFX1 \img_buff_reg[62][5]  ( .D(datain[5]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][5] ) );
  EDFFX1 \img_buff_reg[62][4]  ( .D(datain[4]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][4] ) );
  EDFFX1 \img_buff_reg[62][3]  ( .D(datain[3]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][3] ) );
  EDFFX1 \img_buff_reg[62][2]  ( .D(datain[2]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][2] ) );
  EDFFX1 \img_buff_reg[62][1]  ( .D(datain[1]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][1] ) );
  EDFFX1 \img_buff_reg[62][0]  ( .D(datain[0]), .E(n2355), .CK(clk), .Q(
        \img_buff[62][0] ) );
  EDFFX1 \img_buff_reg[69][7]  ( .D(datain[7]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][7] ) );
  EDFFX1 \img_buff_reg[69][6]  ( .D(datain[6]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][6] ) );
  EDFFX1 \img_buff_reg[69][5]  ( .D(datain[5]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][5] ) );
  EDFFX1 \img_buff_reg[69][4]  ( .D(datain[4]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][4] ) );
  EDFFX1 \img_buff_reg[69][3]  ( .D(datain[3]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][3] ) );
  EDFFX1 \img_buff_reg[69][2]  ( .D(datain[2]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][2] ) );
  EDFFX1 \img_buff_reg[69][1]  ( .D(datain[1]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][1] ) );
  EDFFX1 \img_buff_reg[69][0]  ( .D(datain[0]), .E(n2348), .CK(clk), .Q(
        \img_buff[69][0] ) );
  EDFFX1 \img_buff_reg[72][7]  ( .D(datain[7]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][7] ) );
  EDFFX1 \img_buff_reg[72][6]  ( .D(datain[6]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][6] ) );
  EDFFX1 \img_buff_reg[72][5]  ( .D(datain[5]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][5] ) );
  EDFFX1 \img_buff_reg[72][4]  ( .D(datain[4]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][4] ) );
  EDFFX1 \img_buff_reg[72][3]  ( .D(datain[3]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][3] ) );
  EDFFX1 \img_buff_reg[72][2]  ( .D(datain[2]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][2] ) );
  EDFFX1 \img_buff_reg[72][1]  ( .D(datain[1]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][1] ) );
  EDFFX1 \img_buff_reg[72][0]  ( .D(datain[0]), .E(n2345), .CK(clk), .Q(
        \img_buff[72][0] ) );
  EDFFX1 \img_buff_reg[74][7]  ( .D(datain[7]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][7] ) );
  EDFFX1 \img_buff_reg[74][6]  ( .D(datain[6]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][6] ) );
  EDFFX1 \img_buff_reg[74][5]  ( .D(datain[5]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][5] ) );
  EDFFX1 \img_buff_reg[74][4]  ( .D(datain[4]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][4] ) );
  EDFFX1 \img_buff_reg[74][3]  ( .D(datain[3]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][3] ) );
  EDFFX1 \img_buff_reg[74][2]  ( .D(datain[2]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][2] ) );
  EDFFX1 \img_buff_reg[74][1]  ( .D(datain[1]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][1] ) );
  EDFFX1 \img_buff_reg[74][0]  ( .D(datain[0]), .E(n2343), .CK(clk), .Q(
        \img_buff[74][0] ) );
  EDFFX1 \img_buff_reg[81][7]  ( .D(datain[7]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][7] ) );
  EDFFX1 \img_buff_reg[81][6]  ( .D(datain[6]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][6] ) );
  EDFFX1 \img_buff_reg[81][5]  ( .D(datain[5]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][5] ) );
  EDFFX1 \img_buff_reg[81][4]  ( .D(datain[4]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][4] ) );
  EDFFX1 \img_buff_reg[81][3]  ( .D(datain[3]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][3] ) );
  EDFFX1 \img_buff_reg[81][2]  ( .D(datain[2]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][2] ) );
  EDFFX1 \img_buff_reg[81][1]  ( .D(datain[1]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][1] ) );
  EDFFX1 \img_buff_reg[81][0]  ( .D(datain[0]), .E(n2336), .CK(clk), .Q(
        \img_buff[81][0] ) );
  EDFFX1 \img_buff_reg[89][7]  ( .D(datain[7]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][7] ) );
  EDFFX1 \img_buff_reg[89][6]  ( .D(datain[6]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][6] ) );
  EDFFX1 \img_buff_reg[89][5]  ( .D(datain[5]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][5] ) );
  EDFFX1 \img_buff_reg[89][4]  ( .D(datain[4]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][4] ) );
  EDFFX1 \img_buff_reg[89][3]  ( .D(datain[3]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][3] ) );
  EDFFX1 \img_buff_reg[89][2]  ( .D(datain[2]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][2] ) );
  EDFFX1 \img_buff_reg[89][1]  ( .D(datain[1]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][1] ) );
  EDFFX1 \img_buff_reg[89][0]  ( .D(datain[0]), .E(n2328), .CK(clk), .Q(
        \img_buff[89][0] ) );
  EDFFX1 \img_buff_reg[96][7]  ( .D(datain[7]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][7] ) );
  EDFFX1 \img_buff_reg[96][6]  ( .D(datain[6]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][6] ) );
  EDFFX1 \img_buff_reg[96][5]  ( .D(datain[5]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][5] ) );
  EDFFX1 \img_buff_reg[96][4]  ( .D(datain[4]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][4] ) );
  EDFFX1 \img_buff_reg[96][3]  ( .D(datain[3]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][3] ) );
  EDFFX1 \img_buff_reg[96][2]  ( .D(datain[2]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][2] ) );
  EDFFX1 \img_buff_reg[96][1]  ( .D(datain[1]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][1] ) );
  EDFFX1 \img_buff_reg[96][0]  ( .D(datain[0]), .E(n2321), .CK(clk), .Q(
        \img_buff[96][0] ) );
  EDFFX1 \img_buff_reg[97][7]  ( .D(datain[7]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][7] ) );
  EDFFX1 \img_buff_reg[97][6]  ( .D(datain[6]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][6] ) );
  EDFFX1 \img_buff_reg[97][5]  ( .D(datain[5]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][5] ) );
  EDFFX1 \img_buff_reg[97][4]  ( .D(datain[4]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][4] ) );
  EDFFX1 \img_buff_reg[97][3]  ( .D(datain[3]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][3] ) );
  EDFFX1 \img_buff_reg[97][2]  ( .D(datain[2]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][2] ) );
  EDFFX1 \img_buff_reg[97][1]  ( .D(datain[1]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][1] ) );
  EDFFX1 \img_buff_reg[97][0]  ( .D(datain[0]), .E(n2320), .CK(clk), .Q(
        \img_buff[97][0] ) );
  EDFFX1 \img_buff_reg[101][7]  ( .D(datain[7]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][7] ) );
  EDFFX1 \img_buff_reg[101][6]  ( .D(datain[6]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][6] ) );
  EDFFX1 \img_buff_reg[101][5]  ( .D(datain[5]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][5] ) );
  EDFFX1 \img_buff_reg[101][4]  ( .D(datain[4]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][4] ) );
  EDFFX1 \img_buff_reg[101][3]  ( .D(datain[3]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][3] ) );
  EDFFX1 \img_buff_reg[101][2]  ( .D(datain[2]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][2] ) );
  EDFFX1 \img_buff_reg[101][1]  ( .D(datain[1]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][1] ) );
  EDFFX1 \img_buff_reg[101][0]  ( .D(datain[0]), .E(n2316), .CK(clk), .Q(
        \img_buff[101][0] ) );
  EDFFX1 \img_buff_reg[35][7]  ( .D(datain[7]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][7] ) );
  EDFFX1 \img_buff_reg[35][6]  ( .D(datain[6]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][6] ) );
  EDFFX1 \img_buff_reg[35][5]  ( .D(datain[5]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][5] ) );
  EDFFX1 \img_buff_reg[35][4]  ( .D(datain[4]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][4] ) );
  EDFFX1 \img_buff_reg[35][3]  ( .D(datain[3]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][3] ) );
  EDFFX1 \img_buff_reg[35][2]  ( .D(datain[2]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][2] ) );
  EDFFX1 \img_buff_reg[35][1]  ( .D(datain[1]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][1] ) );
  EDFFX1 \img_buff_reg[35][0]  ( .D(datain[0]), .E(n2382), .CK(clk), .Q(
        \img_buff[35][0] ) );
  EDFFX1 \img_buff_reg[42][7]  ( .D(datain[7]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][7] ) );
  EDFFX1 \img_buff_reg[42][6]  ( .D(datain[6]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][6] ) );
  EDFFX1 \img_buff_reg[42][5]  ( .D(datain[5]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][5] ) );
  EDFFX1 \img_buff_reg[42][4]  ( .D(datain[4]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][4] ) );
  EDFFX1 \img_buff_reg[42][3]  ( .D(datain[3]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][3] ) );
  EDFFX1 \img_buff_reg[42][2]  ( .D(datain[2]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][2] ) );
  EDFFX1 \img_buff_reg[42][1]  ( .D(datain[1]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][1] ) );
  EDFFX1 \img_buff_reg[42][0]  ( .D(datain[0]), .E(n2375), .CK(clk), .Q(
        \img_buff[42][0] ) );
  EDFFX1 \img_buff_reg[43][7]  ( .D(datain[7]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][7] ) );
  EDFFX1 \img_buff_reg[43][6]  ( .D(datain[6]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][6] ) );
  EDFFX1 \img_buff_reg[43][5]  ( .D(datain[5]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][5] ) );
  EDFFX1 \img_buff_reg[43][4]  ( .D(datain[4]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][4] ) );
  EDFFX1 \img_buff_reg[43][3]  ( .D(datain[3]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][3] ) );
  EDFFX1 \img_buff_reg[43][2]  ( .D(datain[2]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][2] ) );
  EDFFX1 \img_buff_reg[43][1]  ( .D(datain[1]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][1] ) );
  EDFFX1 \img_buff_reg[43][0]  ( .D(datain[0]), .E(n2374), .CK(clk), .Q(
        \img_buff[43][0] ) );
  EDFFX1 \img_buff_reg[47][7]  ( .D(datain[7]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][7] ) );
  EDFFX1 \img_buff_reg[47][6]  ( .D(datain[6]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][6] ) );
  EDFFX1 \img_buff_reg[47][5]  ( .D(datain[5]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][5] ) );
  EDFFX1 \img_buff_reg[47][4]  ( .D(datain[4]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][4] ) );
  EDFFX1 \img_buff_reg[47][3]  ( .D(datain[3]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][3] ) );
  EDFFX1 \img_buff_reg[47][2]  ( .D(datain[2]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][2] ) );
  EDFFX1 \img_buff_reg[47][1]  ( .D(datain[1]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][1] ) );
  EDFFX1 \img_buff_reg[47][0]  ( .D(datain[0]), .E(n2370), .CK(clk), .Q(
        \img_buff[47][0] ) );
  EDFFX1 \img_buff_reg[2][7]  ( .D(datain[7]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][7] ) );
  EDFFX1 \img_buff_reg[2][6]  ( .D(datain[6]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][6] ) );
  EDFFX1 \img_buff_reg[2][5]  ( .D(datain[5]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][5] ) );
  EDFFX1 \img_buff_reg[2][4]  ( .D(datain[4]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][4] ) );
  EDFFX1 \img_buff_reg[2][3]  ( .D(datain[3]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][3] ) );
  EDFFX1 \img_buff_reg[2][2]  ( .D(datain[2]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][2] ) );
  EDFFX1 \img_buff_reg[2][1]  ( .D(datain[1]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][1] ) );
  EDFFX1 \img_buff_reg[2][0]  ( .D(datain[0]), .E(n2415), .CK(clk), .Q(
        \img_buff[2][0] ) );
  EDFFX1 \img_buff_reg[7][7]  ( .D(datain[7]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][7] ) );
  EDFFX1 \img_buff_reg[7][6]  ( .D(datain[6]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][6] ) );
  EDFFX1 \img_buff_reg[7][5]  ( .D(datain[5]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][5] ) );
  EDFFX1 \img_buff_reg[7][4]  ( .D(datain[4]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][4] ) );
  EDFFX1 \img_buff_reg[7][3]  ( .D(datain[3]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][3] ) );
  EDFFX1 \img_buff_reg[7][2]  ( .D(datain[2]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][2] ) );
  EDFFX1 \img_buff_reg[7][1]  ( .D(datain[1]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][1] ) );
  EDFFX1 \img_buff_reg[7][0]  ( .D(datain[0]), .E(n2410), .CK(clk), .Q(
        \img_buff[7][0] ) );
  EDFFX1 \img_buff_reg[14][7]  ( .D(datain[7]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][7] ) );
  EDFFX1 \img_buff_reg[14][6]  ( .D(datain[6]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][6] ) );
  EDFFX1 \img_buff_reg[14][5]  ( .D(datain[5]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][5] ) );
  EDFFX1 \img_buff_reg[14][4]  ( .D(datain[4]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][4] ) );
  EDFFX1 \img_buff_reg[14][3]  ( .D(datain[3]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][3] ) );
  EDFFX1 \img_buff_reg[14][2]  ( .D(datain[2]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][2] ) );
  EDFFX1 \img_buff_reg[14][1]  ( .D(datain[1]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][1] ) );
  EDFFX1 \img_buff_reg[14][0]  ( .D(datain[0]), .E(n2403), .CK(clk), .Q(
        \img_buff[14][0] ) );
  EDFFX1 \img_buff_reg[18][7]  ( .D(datain[7]), .E(n2399), .CK(clk), .Q(n2293)
         );
  EDFFX1 \img_buff_reg[18][6]  ( .D(datain[6]), .E(n2399), .CK(clk), .Q(n2259)
         );
  EDFFX1 \img_buff_reg[18][5]  ( .D(datain[5]), .E(n2399), .CK(clk), .Q(n2225)
         );
  EDFFX1 \img_buff_reg[18][4]  ( .D(datain[4]), .E(n2399), .CK(clk), .Q(n2191)
         );
  EDFFX1 \img_buff_reg[18][3]  ( .D(datain[3]), .E(n2399), .CK(clk), .Q(n2157)
         );
  EDFFX1 \img_buff_reg[18][2]  ( .D(datain[2]), .E(n2399), .CK(clk), .Q(n2123)
         );
  EDFFX1 \img_buff_reg[18][1]  ( .D(datain[1]), .E(n2399), .CK(clk), .Q(n2089)
         );
  EDFFX1 \img_buff_reg[18][0]  ( .D(datain[0]), .E(n2399), .CK(clk), .Q(n2055)
         );
  EDFFX1 \img_buff_reg[22][7]  ( .D(datain[7]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][7] ) );
  EDFFX1 \img_buff_reg[22][6]  ( .D(datain[6]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][6] ) );
  EDFFX1 \img_buff_reg[22][5]  ( .D(datain[5]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][5] ) );
  EDFFX1 \img_buff_reg[22][4]  ( .D(datain[4]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][4] ) );
  EDFFX1 \img_buff_reg[22][3]  ( .D(datain[3]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][3] ) );
  EDFFX1 \img_buff_reg[22][2]  ( .D(datain[2]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][2] ) );
  EDFFX1 \img_buff_reg[22][1]  ( .D(datain[1]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][1] ) );
  EDFFX1 \img_buff_reg[22][0]  ( .D(datain[0]), .E(n2395), .CK(clk), .Q(
        \img_buff[22][0] ) );
  EDFFX1 \img_buff_reg[29][7]  ( .D(datain[7]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][7] ) );
  EDFFX1 \img_buff_reg[29][6]  ( .D(datain[6]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][6] ) );
  EDFFX1 \img_buff_reg[29][5]  ( .D(datain[5]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][5] ) );
  EDFFX1 \img_buff_reg[29][4]  ( .D(datain[4]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][4] ) );
  EDFFX1 \img_buff_reg[29][3]  ( .D(datain[3]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][3] ) );
  EDFFX1 \img_buff_reg[29][2]  ( .D(datain[2]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][2] ) );
  EDFFX1 \img_buff_reg[29][1]  ( .D(datain[1]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][1] ) );
  EDFFX1 \img_buff_reg[29][0]  ( .D(datain[0]), .E(n2388), .CK(clk), .Q(
        \img_buff[29][0] ) );
  EDFFX1 \img_buff_reg[49][7]  ( .D(datain[7]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][7] ) );
  EDFFX1 \img_buff_reg[49][6]  ( .D(datain[6]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][6] ) );
  EDFFX1 \img_buff_reg[49][5]  ( .D(datain[5]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][5] ) );
  EDFFX1 \img_buff_reg[49][4]  ( .D(datain[4]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][4] ) );
  EDFFX1 \img_buff_reg[49][3]  ( .D(datain[3]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][3] ) );
  EDFFX1 \img_buff_reg[49][2]  ( .D(datain[2]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][2] ) );
  EDFFX1 \img_buff_reg[49][1]  ( .D(datain[1]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][1] ) );
  EDFFX1 \img_buff_reg[49][0]  ( .D(datain[0]), .E(n2368), .CK(clk), .Q(
        \img_buff[49][0] ) );
  EDFFX1 \img_buff_reg[56][7]  ( .D(datain[7]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][7] ) );
  EDFFX1 \img_buff_reg[56][6]  ( .D(datain[6]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][6] ) );
  EDFFX1 \img_buff_reg[56][5]  ( .D(datain[5]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][5] ) );
  EDFFX1 \img_buff_reg[56][4]  ( .D(datain[4]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][4] ) );
  EDFFX1 \img_buff_reg[56][3]  ( .D(datain[3]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][3] ) );
  EDFFX1 \img_buff_reg[56][2]  ( .D(datain[2]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][2] ) );
  EDFFX1 \img_buff_reg[56][1]  ( .D(datain[1]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][1] ) );
  EDFFX1 \img_buff_reg[56][0]  ( .D(datain[0]), .E(n2361), .CK(clk), .Q(
        \img_buff[56][0] ) );
  EDFFX1 \img_buff_reg[61][7]  ( .D(datain[7]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][7] ) );
  EDFFX1 \img_buff_reg[61][6]  ( .D(datain[6]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][6] ) );
  EDFFX1 \img_buff_reg[61][5]  ( .D(datain[5]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][5] ) );
  EDFFX1 \img_buff_reg[61][4]  ( .D(datain[4]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][4] ) );
  EDFFX1 \img_buff_reg[61][3]  ( .D(datain[3]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][3] ) );
  EDFFX1 \img_buff_reg[61][2]  ( .D(datain[2]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][2] ) );
  EDFFX1 \img_buff_reg[61][1]  ( .D(datain[1]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][1] ) );
  EDFFX1 \img_buff_reg[61][0]  ( .D(datain[0]), .E(n2356), .CK(clk), .Q(
        \img_buff[61][0] ) );
  EDFFX1 \img_buff_reg[68][7]  ( .D(datain[7]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][7] ) );
  EDFFX1 \img_buff_reg[68][6]  ( .D(datain[6]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][6] ) );
  EDFFX1 \img_buff_reg[68][5]  ( .D(datain[5]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][5] ) );
  EDFFX1 \img_buff_reg[68][4]  ( .D(datain[4]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][4] ) );
  EDFFX1 \img_buff_reg[68][3]  ( .D(datain[3]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][3] ) );
  EDFFX1 \img_buff_reg[68][2]  ( .D(datain[2]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][2] ) );
  EDFFX1 \img_buff_reg[68][1]  ( .D(datain[1]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][1] ) );
  EDFFX1 \img_buff_reg[68][0]  ( .D(datain[0]), .E(n2349), .CK(clk), .Q(
        \img_buff[68][0] ) );
  EDFFX1 \img_buff_reg[70][0]  ( .D(datain[0]), .E(n2347), .CK(clk), .Q(n2037)
         );
  EDFFX1 \img_buff_reg[70][7]  ( .D(datain[7]), .E(n2347), .CK(clk), .Q(n2275)
         );
  EDFFX1 \img_buff_reg[70][6]  ( .D(datain[6]), .E(n2347), .CK(clk), .Q(n2241)
         );
  EDFFX1 \img_buff_reg[70][5]  ( .D(datain[5]), .E(n2347), .CK(clk), .Q(n2207)
         );
  EDFFX1 \img_buff_reg[70][4]  ( .D(datain[4]), .E(n2347), .CK(clk), .Q(n2173)
         );
  EDFFX1 \img_buff_reg[70][3]  ( .D(datain[3]), .E(n2347), .CK(clk), .Q(n2139)
         );
  EDFFX1 \img_buff_reg[70][2]  ( .D(datain[2]), .E(n2347), .CK(clk), .Q(n2105)
         );
  EDFFX1 \img_buff_reg[70][1]  ( .D(datain[1]), .E(n2347), .CK(clk), .Q(n2071)
         );
  EDFFX1 \img_buff_reg[76][7]  ( .D(datain[7]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][7] ) );
  EDFFX1 \img_buff_reg[76][6]  ( .D(datain[6]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][6] ) );
  EDFFX1 \img_buff_reg[76][5]  ( .D(datain[5]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][5] ) );
  EDFFX1 \img_buff_reg[76][4]  ( .D(datain[4]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][4] ) );
  EDFFX1 \img_buff_reg[76][3]  ( .D(datain[3]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][3] ) );
  EDFFX1 \img_buff_reg[76][2]  ( .D(datain[2]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][2] ) );
  EDFFX1 \img_buff_reg[76][1]  ( .D(datain[1]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][1] ) );
  EDFFX1 \img_buff_reg[76][0]  ( .D(datain[0]), .E(n2341), .CK(clk), .Q(
        \img_buff[76][0] ) );
  EDFFX1 \img_buff_reg[83][5]  ( .D(datain[5]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][5] ) );
  EDFFX1 \img_buff_reg[83][4]  ( .D(datain[4]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][4] ) );
  EDFFX1 \img_buff_reg[83][3]  ( .D(datain[3]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][3] ) );
  EDFFX1 \img_buff_reg[83][2]  ( .D(datain[2]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][2] ) );
  EDFFX1 \img_buff_reg[83][1]  ( .D(datain[1]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][1] ) );
  EDFFX1 \img_buff_reg[83][0]  ( .D(datain[0]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][0] ) );
  EDFFX1 \img_buff_reg[83][7]  ( .D(datain[7]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][7] ) );
  EDFFX1 \img_buff_reg[83][6]  ( .D(datain[6]), .E(n2334), .CK(clk), .Q(
        \img_buff[83][6] ) );
  EDFFX1 \img_buff_reg[88][7]  ( .D(datain[7]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][7] ) );
  EDFFX1 \img_buff_reg[88][6]  ( .D(datain[6]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][6] ) );
  EDFFX1 \img_buff_reg[88][5]  ( .D(datain[5]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][5] ) );
  EDFFX1 \img_buff_reg[88][4]  ( .D(datain[4]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][4] ) );
  EDFFX1 \img_buff_reg[88][3]  ( .D(datain[3]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][3] ) );
  EDFFX1 \img_buff_reg[88][2]  ( .D(datain[2]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][2] ) );
  EDFFX1 \img_buff_reg[88][1]  ( .D(datain[1]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][1] ) );
  EDFFX1 \img_buff_reg[88][0]  ( .D(datain[0]), .E(n2329), .CK(clk), .Q(
        \img_buff[88][0] ) );
  EDFFX1 \img_buff_reg[95][2]  ( .D(datain[2]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][2] ) );
  EDFFX1 \img_buff_reg[95][1]  ( .D(datain[1]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][1] ) );
  EDFFX1 \img_buff_reg[95][0]  ( .D(datain[0]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][0] ) );
  EDFFX1 \img_buff_reg[95][7]  ( .D(datain[7]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][7] ) );
  EDFFX1 \img_buff_reg[95][6]  ( .D(datain[6]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][6] ) );
  EDFFX1 \img_buff_reg[95][5]  ( .D(datain[5]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][5] ) );
  EDFFX1 \img_buff_reg[95][4]  ( .D(datain[4]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][4] ) );
  EDFFX1 \img_buff_reg[95][3]  ( .D(datain[3]), .E(n2322), .CK(clk), .Q(
        \img_buff[95][3] ) );
  EDFFX1 \img_buff_reg[99][7]  ( .D(datain[7]), .E(n2318), .CK(clk), .Q(n2285)
         );
  EDFFX1 \img_buff_reg[99][6]  ( .D(datain[6]), .E(n2318), .CK(clk), .Q(n2251)
         );
  EDFFX1 \img_buff_reg[99][5]  ( .D(datain[5]), .E(n2318), .CK(clk), .Q(n2217)
         );
  EDFFX1 \img_buff_reg[99][4]  ( .D(datain[4]), .E(n2318), .CK(clk), .Q(n2183)
         );
  EDFFX1 \img_buff_reg[99][3]  ( .D(datain[3]), .E(n2318), .CK(clk), .Q(n2149)
         );
  EDFFX1 \img_buff_reg[99][2]  ( .D(datain[2]), .E(n2318), .CK(clk), .Q(n2115)
         );
  EDFFX1 \img_buff_reg[99][1]  ( .D(datain[1]), .E(n2318), .CK(clk), .Q(n2081)
         );
  EDFFX1 \img_buff_reg[99][0]  ( .D(datain[0]), .E(n2318), .CK(clk), .Q(n2047)
         );
  EDFFX1 \img_buff_reg[103][7]  ( .D(datain[7]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][7] ) );
  EDFFX1 \img_buff_reg[103][6]  ( .D(datain[6]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][6] ) );
  EDFFX1 \img_buff_reg[103][5]  ( .D(datain[5]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][5] ) );
  EDFFX1 \img_buff_reg[103][4]  ( .D(datain[4]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][4] ) );
  EDFFX1 \img_buff_reg[103][3]  ( .D(datain[3]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][3] ) );
  EDFFX1 \img_buff_reg[103][2]  ( .D(datain[2]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][2] ) );
  EDFFX1 \img_buff_reg[103][1]  ( .D(datain[1]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][1] ) );
  EDFFX1 \img_buff_reg[103][0]  ( .D(datain[0]), .E(n2314), .CK(clk), .Q(
        \img_buff[103][0] ) );
  EDFFX1 \img_buff_reg[34][7]  ( .D(datain[7]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][7] ) );
  EDFFX1 \img_buff_reg[34][6]  ( .D(datain[6]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][6] ) );
  EDFFX1 \img_buff_reg[34][5]  ( .D(datain[5]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][5] ) );
  EDFFX1 \img_buff_reg[34][4]  ( .D(datain[4]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][4] ) );
  EDFFX1 \img_buff_reg[34][3]  ( .D(datain[3]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][3] ) );
  EDFFX1 \img_buff_reg[34][2]  ( .D(datain[2]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][2] ) );
  EDFFX1 \img_buff_reg[34][1]  ( .D(datain[1]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][1] ) );
  EDFFX1 \img_buff_reg[34][0]  ( .D(datain[0]), .E(n2383), .CK(clk), .Q(
        \img_buff[34][0] ) );
  EDFFX1 \img_buff_reg[41][7]  ( .D(datain[7]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][7] ) );
  EDFFX1 \img_buff_reg[41][6]  ( .D(datain[6]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][6] ) );
  EDFFX1 \img_buff_reg[41][5]  ( .D(datain[5]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][5] ) );
  EDFFX1 \img_buff_reg[41][4]  ( .D(datain[4]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][4] ) );
  EDFFX1 \img_buff_reg[41][3]  ( .D(datain[3]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][3] ) );
  EDFFX1 \img_buff_reg[41][2]  ( .D(datain[2]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][2] ) );
  EDFFX1 \img_buff_reg[41][1]  ( .D(datain[1]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][1] ) );
  EDFFX1 \img_buff_reg[41][0]  ( .D(datain[0]), .E(n2376), .CK(clk), .Q(
        \img_buff[41][0] ) );
  EDFFX1 \img_buff_reg[45][7]  ( .D(datain[7]), .E(n2372), .CK(clk), .Q(n2301)
         );
  EDFFX1 \img_buff_reg[45][6]  ( .D(datain[6]), .E(n2372), .CK(clk), .Q(n2267)
         );
  EDFFX1 \img_buff_reg[45][5]  ( .D(datain[5]), .E(n2372), .CK(clk), .Q(n2233)
         );
  EDFFX1 \img_buff_reg[45][4]  ( .D(datain[4]), .E(n2372), .CK(clk), .Q(n2199)
         );
  EDFFX1 \img_buff_reg[45][3]  ( .D(datain[3]), .E(n2372), .CK(clk), .Q(n2165)
         );
  EDFFX1 \img_buff_reg[45][2]  ( .D(datain[2]), .E(n2372), .CK(clk), .Q(n2131)
         );
  EDFFX1 \img_buff_reg[45][1]  ( .D(datain[1]), .E(n2372), .CK(clk), .Q(n2097)
         );
  EDFFX1 \img_buff_reg[45][0]  ( .D(datain[0]), .E(n2372), .CK(clk), .Q(n2063)
         );
  EDFFX1 \img_buff_reg[6][7]  ( .D(datain[7]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][7] ) );
  EDFFX1 \img_buff_reg[6][6]  ( .D(datain[6]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][6] ) );
  EDFFX1 \img_buff_reg[6][5]  ( .D(datain[5]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][5] ) );
  EDFFX1 \img_buff_reg[6][4]  ( .D(datain[4]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][4] ) );
  EDFFX1 \img_buff_reg[6][3]  ( .D(datain[3]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][3] ) );
  EDFFX1 \img_buff_reg[6][2]  ( .D(datain[2]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][2] ) );
  EDFFX1 \img_buff_reg[6][1]  ( .D(datain[1]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][1] ) );
  EDFFX1 \img_buff_reg[6][0]  ( .D(datain[0]), .E(n2411), .CK(clk), .Q(
        \img_buff[6][0] ) );
  EDFFX1 \img_buff_reg[13][7]  ( .D(datain[7]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][7] ) );
  EDFFX1 \img_buff_reg[13][6]  ( .D(datain[6]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][6] ) );
  EDFFX1 \img_buff_reg[13][5]  ( .D(datain[5]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][5] ) );
  EDFFX1 \img_buff_reg[13][4]  ( .D(datain[4]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][4] ) );
  EDFFX1 \img_buff_reg[13][3]  ( .D(datain[3]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][3] ) );
  EDFFX1 \img_buff_reg[13][2]  ( .D(datain[2]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][2] ) );
  EDFFX1 \img_buff_reg[13][1]  ( .D(datain[1]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][1] ) );
  EDFFX1 \img_buff_reg[13][0]  ( .D(datain[0]), .E(n2404), .CK(clk), .Q(
        \img_buff[13][0] ) );
  EDFFX1 \img_buff_reg[17][7]  ( .D(datain[7]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][7] ) );
  EDFFX1 \img_buff_reg[17][6]  ( .D(datain[6]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][6] ) );
  EDFFX1 \img_buff_reg[17][5]  ( .D(datain[5]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][5] ) );
  EDFFX1 \img_buff_reg[17][4]  ( .D(datain[4]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][4] ) );
  EDFFX1 \img_buff_reg[17][3]  ( .D(datain[3]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][3] ) );
  EDFFX1 \img_buff_reg[17][2]  ( .D(datain[2]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][2] ) );
  EDFFX1 \img_buff_reg[17][1]  ( .D(datain[1]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][1] ) );
  EDFFX1 \img_buff_reg[17][0]  ( .D(datain[0]), .E(n2400), .CK(clk), .Q(
        \img_buff[17][0] ) );
  EDFFX1 \img_buff_reg[60][7]  ( .D(datain[7]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][7] ) );
  EDFFX1 \img_buff_reg[60][6]  ( .D(datain[6]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][6] ) );
  EDFFX1 \img_buff_reg[60][5]  ( .D(datain[5]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][5] ) );
  EDFFX1 \img_buff_reg[60][4]  ( .D(datain[4]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][4] ) );
  EDFFX1 \img_buff_reg[60][3]  ( .D(datain[3]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][3] ) );
  EDFFX1 \img_buff_reg[60][2]  ( .D(datain[2]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][2] ) );
  EDFFX1 \img_buff_reg[60][1]  ( .D(datain[1]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][1] ) );
  EDFFX1 \img_buff_reg[60][0]  ( .D(datain[0]), .E(n2357), .CK(clk), .Q(
        \img_buff[60][0] ) );
  EDFFX1 \img_buff_reg[67][7]  ( .D(datain[7]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][7] ) );
  EDFFX1 \img_buff_reg[67][6]  ( .D(datain[6]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][6] ) );
  EDFFX1 \img_buff_reg[67][5]  ( .D(datain[5]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][5] ) );
  EDFFX1 \img_buff_reg[67][4]  ( .D(datain[4]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][4] ) );
  EDFFX1 \img_buff_reg[67][3]  ( .D(datain[3]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][3] ) );
  EDFFX1 \img_buff_reg[67][2]  ( .D(datain[2]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][2] ) );
  EDFFX1 \img_buff_reg[67][1]  ( .D(datain[1]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][1] ) );
  EDFFX1 \img_buff_reg[67][0]  ( .D(datain[0]), .E(n2350), .CK(clk), .Q(
        \img_buff[67][0] ) );
  EDFFX1 \img_buff_reg[73][7]  ( .D(datain[7]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][7] ) );
  EDFFX1 \img_buff_reg[73][6]  ( .D(datain[6]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][6] ) );
  EDFFX1 \img_buff_reg[73][5]  ( .D(datain[5]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][5] ) );
  EDFFX1 \img_buff_reg[73][4]  ( .D(datain[4]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][4] ) );
  EDFFX1 \img_buff_reg[73][3]  ( .D(datain[3]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][3] ) );
  EDFFX1 \img_buff_reg[73][2]  ( .D(datain[2]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][2] ) );
  EDFFX1 \img_buff_reg[73][1]  ( .D(datain[1]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][1] ) );
  EDFFX1 \img_buff_reg[73][0]  ( .D(datain[0]), .E(n2344), .CK(clk), .Q(
        \img_buff[73][0] ) );
  EDFFX1 \img_buff_reg[87][7]  ( .D(datain[7]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][7] ) );
  EDFFX1 \img_buff_reg[87][6]  ( .D(datain[6]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][6] ) );
  EDFFX1 \img_buff_reg[87][5]  ( .D(datain[5]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][5] ) );
  EDFFX1 \img_buff_reg[87][4]  ( .D(datain[4]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][4] ) );
  EDFFX1 \img_buff_reg[87][3]  ( .D(datain[3]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][3] ) );
  EDFFX1 \img_buff_reg[87][2]  ( .D(datain[2]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][2] ) );
  EDFFX1 \img_buff_reg[87][1]  ( .D(datain[1]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][1] ) );
  EDFFX1 \img_buff_reg[87][0]  ( .D(datain[0]), .E(n2330), .CK(clk), .Q(
        \img_buff[87][0] ) );
  EDFFX1 \img_buff_reg[94][7]  ( .D(datain[7]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][7] ) );
  EDFFX1 \img_buff_reg[94][6]  ( .D(datain[6]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][6] ) );
  EDFFX1 \img_buff_reg[94][5]  ( .D(datain[5]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][5] ) );
  EDFFX1 \img_buff_reg[94][4]  ( .D(datain[4]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][4] ) );
  EDFFX1 \img_buff_reg[94][3]  ( .D(datain[3]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][3] ) );
  EDFFX1 \img_buff_reg[94][2]  ( .D(datain[2]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][2] ) );
  EDFFX1 \img_buff_reg[94][1]  ( .D(datain[1]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][1] ) );
  EDFFX1 \img_buff_reg[94][0]  ( .D(datain[0]), .E(n2323), .CK(clk), .Q(
        \img_buff[94][0] ) );
  EDFFX1 \img_buff_reg[98][7]  ( .D(datain[7]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][7] ) );
  EDFFX1 \img_buff_reg[98][6]  ( .D(datain[6]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][6] ) );
  EDFFX1 \img_buff_reg[98][5]  ( .D(datain[5]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][5] ) );
  EDFFX1 \img_buff_reg[98][4]  ( .D(datain[4]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][4] ) );
  EDFFX1 \img_buff_reg[98][3]  ( .D(datain[3]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][3] ) );
  EDFFX1 \img_buff_reg[98][2]  ( .D(datain[2]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][2] ) );
  EDFFX1 \img_buff_reg[98][1]  ( .D(datain[1]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][1] ) );
  EDFFX1 \img_buff_reg[98][0]  ( .D(datain[0]), .E(n2319), .CK(clk), .Q(
        \img_buff[98][0] ) );
  EDFFX1 \img_buff_reg[33][1]  ( .D(datain[1]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][1] ) );
  EDFFX1 \img_buff_reg[33][0]  ( .D(datain[0]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][0] ) );
  EDFFX1 \img_buff_reg[33][7]  ( .D(datain[7]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][7] ) );
  EDFFX1 \img_buff_reg[33][6]  ( .D(datain[6]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][6] ) );
  EDFFX1 \img_buff_reg[33][5]  ( .D(datain[5]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][5] ) );
  EDFFX1 \img_buff_reg[33][4]  ( .D(datain[4]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][4] ) );
  EDFFX1 \img_buff_reg[33][3]  ( .D(datain[3]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][3] ) );
  EDFFX1 \img_buff_reg[33][2]  ( .D(datain[2]), .E(n2384), .CK(clk), .Q(
        \img_buff[33][2] ) );
  EDFFX1 \img_buff_reg[40][7]  ( .D(datain[7]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][7] ) );
  EDFFX1 \img_buff_reg[40][6]  ( .D(datain[6]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][6] ) );
  EDFFX1 \img_buff_reg[40][5]  ( .D(datain[5]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][5] ) );
  EDFFX1 \img_buff_reg[40][4]  ( .D(datain[4]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][4] ) );
  EDFFX1 \img_buff_reg[40][3]  ( .D(datain[3]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][3] ) );
  EDFFX1 \img_buff_reg[40][2]  ( .D(datain[2]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][2] ) );
  EDFFX1 \img_buff_reg[40][1]  ( .D(datain[1]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][1] ) );
  EDFFX1 \img_buff_reg[40][0]  ( .D(datain[0]), .E(n2377), .CK(clk), .Q(
        \img_buff[40][0] ) );
  EDFFX1 \img_buff_reg[44][7]  ( .D(datain[7]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][7] ) );
  EDFFX1 \img_buff_reg[44][6]  ( .D(datain[6]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][6] ) );
  EDFFX1 \img_buff_reg[44][5]  ( .D(datain[5]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][5] ) );
  EDFFX1 \img_buff_reg[44][4]  ( .D(datain[4]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][4] ) );
  EDFFX1 \img_buff_reg[44][3]  ( .D(datain[3]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][3] ) );
  EDFFX1 \img_buff_reg[44][2]  ( .D(datain[2]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][2] ) );
  EDFFX1 \img_buff_reg[44][1]  ( .D(datain[1]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][1] ) );
  EDFFX1 \img_buff_reg[44][0]  ( .D(datain[0]), .E(n2373), .CK(clk), .Q(
        \img_buff[44][0] ) );
  DFFRXL output_valid_reg ( .D(n1267), .CK(clk), .RN(n2309), .Q(output_valid), 
        .QN(n2303) );
  DFFRXL busy_reg ( .D(n1266), .CK(clk), .RN(n2309), .Q(busy), .QN(n2302) );
  DFFRXL \img_counter_reg[7]  ( .D(n1278), .CK(clk), .RN(n2309), .Q(
        img_counter[7]), .QN(n224) );
  DFFRXL \dataout_reg[0]  ( .D(n1254), .CK(clk), .RN(n2309), .Q(dataout[0]) );
  DFFRXL \dataout_reg[1]  ( .D(n1255), .CK(clk), .RN(n2309), .Q(dataout[1]) );
  DFFRXL \dataout_reg[2]  ( .D(n1256), .CK(clk), .RN(n2309), .Q(dataout[2]) );
  DFFRXL \dataout_reg[3]  ( .D(n1257), .CK(clk), .RN(n2309), .Q(dataout[3]) );
  DFFRXL \dataout_reg[4]  ( .D(n1258), .CK(clk), .RN(n2309), .Q(dataout[4]) );
  DFFRXL \dataout_reg[5]  ( .D(n1259), .CK(clk), .RN(n2309), .Q(dataout[5]) );
  DFFRXL \dataout_reg[6]  ( .D(n1260), .CK(clk), .RN(n2309), .Q(dataout[6]) );
  DFFRXL \dataout_reg[7]  ( .D(n1261), .CK(clk), .RN(n2309), .Q(dataout[7]) );
  DFFRXL \L_reg[0]  ( .D(n1265), .CK(clk), .RN(n2309), .Q(n2304), .QN(n1286)
         );
  DFFRXL \img_counter_reg[5]  ( .D(n1271), .CK(clk), .RN(n2309), .Q(
        img_counter[5]), .QN(n226) );
  DFFRXL \img_counter_reg[6]  ( .D(n1270), .CK(clk), .RN(n2309), .Q(
        img_counter[6]), .QN(n225) );
  DFFRXL \img_counter_reg[1]  ( .D(n1275), .CK(clk), .RN(n2309), .Q(
        img_counter[1]), .QN(n230) );
  DFFRXL \img_counter_reg[2]  ( .D(n1274), .CK(clk), .RN(n2309), .Q(
        img_counter[2]), .QN(n229) );
  DFFRXL \img_counter_reg[3]  ( .D(n1273), .CK(clk), .RN(n2309), .Q(
        img_counter[3]), .QN(n228) );
  DFFRXL \img_counter_reg[4]  ( .D(n1272), .CK(clk), .RN(n2309), .Q(
        img_counter[4]), .QN(n227) );
  DFFRXL \img_counter_reg[0]  ( .D(n1276), .CK(clk), .RN(n2309), .Q(
        img_counter[0]), .QN(n231) );
  XOR3X1 \r594/U1_6  ( .A(\U3/U15/Z_5 ), .B(\U3/U15/Z_6 ), .C(\r594/carry[6] ), 
        .Y(N1003) );
  XOR3X1 \r481/U1_6  ( .A(\U3/U16/Z_6 ), .B(N1003), .C(\r481/carry[6] ), .Y(
        out_pos[6]) );
  ADDFXL \r481/U1_5  ( .A(\U3/U16/Z_5 ), .B(N1002), .CI(\r481/carry[5] ), .CO(
        \r481/carry[6] ), .S(out_pos[5]) );
  ADDFXL \r481/U1_4  ( .A(\U3/U16/Z_4 ), .B(N1001), .CI(\r481/carry[4] ), .CO(
        \r481/carry[5] ), .S(out_pos[4]) );
  ADDFXL \r597/U1_2  ( .A(\U3/U10/Z_2 ), .B(\U3/U11/Z_2 ), .CI(\r597/carry[2] ), .CO(\r597/carry[3] ), .S(N983) );
  ADDFXL \r597/U1_1  ( .A(\U3/U10/Z_1 ), .B(\U3/U11/Z_1 ), .CI(\r597/carry[1] ), .CO(\r597/carry[2] ), .S(N982) );
  ADDFXL \r597/U1_3  ( .A(\U3/U10/Z_3 ), .B(\U3/U11/Z_3 ), .CI(\r597/carry[3] ), .CO(\r597/carry[4] ), .S(N984) );
  ADDFXL \r596/U2_2  ( .A(N983), .B(n2306), .CI(\r596/carry[2] ), .CO(
        \r596/carry[3] ), .S(N987) );
  ADDFXL \r596/U2_1  ( .A(N982), .B(n2308), .CI(\r596/carry[1] ), .CO(
        \r596/carry[2] ), .S(out_pos[1]) );
  ADDFXL \r481/U1_3  ( .A(N988), .B(N1000), .CI(\r481/carry[3] ), .CO(
        \r481/carry[4] ), .S(out_pos[3]) );
  ADDFXL \r594/U1_5  ( .A(\U3/U15/Z_4 ), .B(\U3/U15/Z_5 ), .CI(\r594/carry[5] ), .CO(\r594/carry[6] ), .S(N1002) );
  ADDFXL \r594/U1_4  ( .A(\U3/U15/Z_3 ), .B(\U3/U15/Z_4 ), .CI(\r594/carry[4] ), .CO(\r594/carry[5] ), .S(N1001) );
  ADDFXL \r596/U2_3  ( .A(N984), .B(n2305), .CI(\r596/carry[3] ), .CO(
        \r596/carry[4] ), .S(N988) );
  INVX3 U1008 ( .A(reset), .Y(n2309) );
  CLKINVX1 U1009 ( .A(N987), .Y(n1296) );
  NOR2X1 U1010 ( .A(n1287), .B(n2305), .Y(N966) );
  NAND2BX1 U1011 ( .AN(n1300), .B(\U3/U13/Z_2 ), .Y(n1287) );
  XNOR2X1 U1012 ( .A(\U3/U11/Z_0 ), .B(n1291), .Y(N981) );
  XNOR2X1 U1013 ( .A(N999), .B(n1296), .Y(out_pos[2]) );
  XNOR2X1 U1014 ( .A(n2307), .B(N981), .Y(out_pos[0]) );
  CLKINVX1 U1015 ( .A(N999), .Y(n1297) );
  OR2X1 U1016 ( .A(\U3/U12/Z_4 ), .B(\r596/carry[4] ), .Y(\r596/carry[5] ) );
  CLKINVX1 U1017 ( .A(n2307), .Y(n1294) );
  CLKINVX1 U1018 ( .A(\U3/U11/Z_0 ), .Y(n1299) );
  CLKINVX1 U1019 ( .A(\U3/U12/Z_5 ), .Y(n1292) );
  NOR2X1 U1020 ( .A(n1297), .B(n1298), .Y(\r594/carry[4] ) );
  CLKINVX1 U1021 ( .A(\U3/U15/Z_3 ), .Y(n1298) );
  NOR2X1 U1022 ( .A(n1296), .B(n1297), .Y(\r481/carry[3] ) );
  XNOR2X1 U1023 ( .A(\U3/U15/Z_3 ), .B(n1297), .Y(N1000) );
  NAND2X1 U1024 ( .A(n1294), .B(n1295), .Y(\r596/carry[1] ) );
  CLKINVX1 U1025 ( .A(N981), .Y(n1295) );
  CLKINVX1 U1026 ( .A(\r597/carry[4] ), .Y(n1300) );
  NOR2X1 U1027 ( .A(n1288), .B(n1290), .Y(\U3/U12/Z_4 ) );
  XOR2X1 U1028 ( .A(\U3/U13/Z_2 ), .B(n1300), .Y(n1288) );
  NOR2X1 U1029 ( .A(n1289), .B(n1290), .Y(\U3/U12/Z_5 ) );
  XOR2X1 U1030 ( .A(\U3/U13/Z_3 ), .B(n1287), .Y(n1289) );
  XNOR2X1 U1031 ( .A(\U3/U12/Z_6 ), .B(\r596/carry[6] ), .Y(N973) );
  NAND2X1 U1032 ( .A(n1292), .B(n1293), .Y(\r596/carry[6] ) );
  CLKINVX1 U1033 ( .A(\r596/carry[5] ), .Y(n1293) );
  OR2X1 U1034 ( .A(n432), .B(n1286), .Y(n1291) );
  NOR2X1 U1035 ( .A(n1291), .B(n1299), .Y(\r597/carry[1] ) );
  XNOR2X1 U1036 ( .A(\U3/U12/Z_4 ), .B(\r596/carry[4] ), .Y(N971) );
  XNOR2X1 U1037 ( .A(\U3/U12/Z_5 ), .B(\r596/carry[5] ), .Y(N972) );
  NOR2X1 U1038 ( .A(img_counter[1]), .B(n1290), .Y(n2308) );
  OAI2BB1X1 U1039 ( .A0N(n1284), .A1N(n1301), .B0(n1302), .Y(next_state) );
  NOR2X1 U1040 ( .A(n1303), .B(n1304), .Y(n2311) );
  NOR2X1 U1041 ( .A(n1303), .B(n1305), .Y(n2312) );
  NOR2X1 U1042 ( .A(n1303), .B(n1306), .Y(n2313) );
  NOR2X1 U1043 ( .A(n1303), .B(n1307), .Y(n2314) );
  NOR2X1 U1044 ( .A(n1303), .B(n1308), .Y(n2315) );
  NOR2X1 U1045 ( .A(n1303), .B(n1309), .Y(n2316) );
  NOR2X1 U1046 ( .A(n1303), .B(n1310), .Y(n2317) );
  NOR2X1 U1047 ( .A(n1311), .B(n1303), .Y(n2318) );
  NOR2X1 U1048 ( .A(n1303), .B(n1312), .Y(n2319) );
  NOR2X1 U1049 ( .A(n1303), .B(n1313), .Y(n2320) );
  NOR2X1 U1050 ( .A(n1303), .B(n1314), .Y(n2321) );
  NAND3X1 U1051 ( .A(img_counter[6]), .B(img_counter[5]), .C(n1315), .Y(n1303)
         );
  NOR2X1 U1052 ( .A(n1316), .B(n1317), .Y(n2322) );
  NOR2X1 U1053 ( .A(n1316), .B(n1318), .Y(n2323) );
  NOR2X1 U1054 ( .A(n1316), .B(n1319), .Y(n2324) );
  NOR2X1 U1055 ( .A(n1316), .B(n1320), .Y(n2325) );
  NOR2X1 U1056 ( .A(n1321), .B(n1316), .Y(n2326) );
  NOR2X1 U1057 ( .A(n1304), .B(n1316), .Y(n2327) );
  NOR2X1 U1058 ( .A(n1305), .B(n1316), .Y(n2328) );
  NOR2X1 U1059 ( .A(n1306), .B(n1316), .Y(n2329) );
  NOR2X1 U1060 ( .A(n1307), .B(n1316), .Y(n2330) );
  NOR2X1 U1061 ( .A(n1308), .B(n1316), .Y(n2331) );
  NOR2X1 U1062 ( .A(n1309), .B(n1316), .Y(n2332) );
  NOR2X1 U1063 ( .A(n1310), .B(n1316), .Y(n2333) );
  NOR2X1 U1064 ( .A(n1311), .B(n1316), .Y(n2334) );
  NOR2X1 U1065 ( .A(n1312), .B(n1316), .Y(n2335) );
  NOR2X1 U1066 ( .A(n1313), .B(n1316), .Y(n2336) );
  NOR2X1 U1067 ( .A(n1314), .B(n1316), .Y(n2337) );
  NAND2X1 U1068 ( .A(n1322), .B(img_counter[6]), .Y(n1316) );
  NOR2X1 U1069 ( .A(n1317), .B(n1323), .Y(n2338) );
  NOR2X1 U1070 ( .A(n1318), .B(n1323), .Y(n2339) );
  NOR2X1 U1071 ( .A(n1319), .B(n1323), .Y(n2340) );
  NOR2X1 U1072 ( .A(n1320), .B(n1323), .Y(n2341) );
  NOR2X1 U1073 ( .A(n1321), .B(n1323), .Y(n2342) );
  NOR2X1 U1074 ( .A(n1304), .B(n1323), .Y(n2343) );
  NOR2X1 U1075 ( .A(n1305), .B(n1323), .Y(n2344) );
  NOR2X1 U1076 ( .A(n1306), .B(n1323), .Y(n2345) );
  NOR2X1 U1077 ( .A(n1307), .B(n1323), .Y(n2346) );
  NOR2X1 U1078 ( .A(n1308), .B(n1323), .Y(n2347) );
  NOR2X1 U1079 ( .A(n1309), .B(n1323), .Y(n2348) );
  NOR2X1 U1080 ( .A(n1310), .B(n1323), .Y(n2349) );
  NOR2X1 U1081 ( .A(n1311), .B(n1323), .Y(n2350) );
  NOR2X1 U1082 ( .A(n1312), .B(n1323), .Y(n2351) );
  NOR2X1 U1083 ( .A(n1313), .B(n1323), .Y(n2352) );
  NOR2X1 U1084 ( .A(n1314), .B(n1323), .Y(n2353) );
  NAND3X1 U1085 ( .A(n1315), .B(img_counter[6]), .C(n226), .Y(n1323) );
  NOR2X1 U1086 ( .A(n1317), .B(n1324), .Y(n2354) );
  NOR2X1 U1087 ( .A(n1318), .B(n1324), .Y(n2355) );
  NOR2X1 U1088 ( .A(n1319), .B(n1324), .Y(n2356) );
  NOR2X1 U1089 ( .A(n1320), .B(n1324), .Y(n2357) );
  NOR2X1 U1090 ( .A(n1321), .B(n1324), .Y(n2358) );
  NOR2X1 U1091 ( .A(n1304), .B(n1324), .Y(n2359) );
  NOR2X1 U1092 ( .A(n1305), .B(n1324), .Y(n2360) );
  NOR2X1 U1093 ( .A(n1306), .B(n1324), .Y(n2361) );
  NOR2X1 U1094 ( .A(n1307), .B(n1324), .Y(n2362) );
  NOR2X1 U1095 ( .A(n1308), .B(n1324), .Y(n2363) );
  NOR2X1 U1096 ( .A(n1309), .B(n1324), .Y(n2364) );
  NOR2X1 U1097 ( .A(n1310), .B(n1324), .Y(n2365) );
  NOR2X1 U1098 ( .A(n1311), .B(n1324), .Y(n2366) );
  NOR2X1 U1099 ( .A(n1312), .B(n1324), .Y(n2367) );
  NOR2X1 U1100 ( .A(n1313), .B(n1324), .Y(n2368) );
  NOR2X1 U1101 ( .A(n1314), .B(n1324), .Y(n2369) );
  NAND4X1 U1102 ( .A(n1325), .B(n225), .C(img_counter[5]), .D(img_counter[4]), 
        .Y(n1324) );
  NOR2X1 U1103 ( .A(n1317), .B(n1326), .Y(n2370) );
  NOR2X1 U1104 ( .A(n1318), .B(n1326), .Y(n2371) );
  NOR2X1 U1105 ( .A(n1319), .B(n1326), .Y(n2372) );
  NOR2X1 U1106 ( .A(n1320), .B(n1326), .Y(n2373) );
  NOR2X1 U1107 ( .A(n1321), .B(n1326), .Y(n2374) );
  NOR2X1 U1108 ( .A(n1304), .B(n1326), .Y(n2375) );
  NOR2X1 U1109 ( .A(n1305), .B(n1326), .Y(n2376) );
  NOR2X1 U1110 ( .A(n1306), .B(n1326), .Y(n2377) );
  NOR2X1 U1111 ( .A(n1307), .B(n1326), .Y(n2378) );
  NOR2X1 U1112 ( .A(n1308), .B(n1326), .Y(n2379) );
  NOR2X1 U1113 ( .A(n1309), .B(n1326), .Y(n2380) );
  NOR2X1 U1114 ( .A(n1310), .B(n1326), .Y(n2381) );
  NOR2X1 U1115 ( .A(n1311), .B(n1326), .Y(n2382) );
  NOR2X1 U1116 ( .A(n1312), .B(n1326), .Y(n2383) );
  NOR2X1 U1117 ( .A(n1313), .B(n1326), .Y(n2384) );
  NOR2X1 U1118 ( .A(n1314), .B(n1326), .Y(n2385) );
  NAND3X1 U1119 ( .A(n225), .B(img_counter[5]), .C(n1315), .Y(n1326) );
  NOR2X1 U1120 ( .A(n1317), .B(n1327), .Y(n2386) );
  NOR2X1 U1121 ( .A(n1318), .B(n1327), .Y(n2387) );
  NOR2X1 U1122 ( .A(n1319), .B(n1327), .Y(n2388) );
  NOR2X1 U1123 ( .A(n1320), .B(n1327), .Y(n2389) );
  NOR2X1 U1124 ( .A(n1321), .B(n1327), .Y(n2390) );
  NOR2X1 U1125 ( .A(n1304), .B(n1327), .Y(n2391) );
  NOR2X1 U1126 ( .A(n1305), .B(n1327), .Y(n2392) );
  NOR2X1 U1127 ( .A(n1306), .B(n1327), .Y(n2393) );
  NOR2X1 U1128 ( .A(n1307), .B(n1327), .Y(n2394) );
  NOR2X1 U1129 ( .A(n1308), .B(n1327), .Y(n2395) );
  NOR2X1 U1130 ( .A(n1309), .B(n1327), .Y(n2396) );
  NOR2X1 U1131 ( .A(n1310), .B(n1327), .Y(n2397) );
  NOR2X1 U1132 ( .A(n1311), .B(n1327), .Y(n2398) );
  NOR2X1 U1133 ( .A(n1312), .B(n1327), .Y(n2399) );
  NOR2X1 U1134 ( .A(n1313), .B(n1327), .Y(n2400) );
  NOR2X1 U1135 ( .A(n1314), .B(n1327), .Y(n2401) );
  NAND2X1 U1136 ( .A(n1322), .B(n225), .Y(n1327) );
  NOR3BXL U1137 ( .AN(n1325), .B(n227), .C(img_counter[5]), .Y(n1322) );
  NOR2X1 U1138 ( .A(n1317), .B(n1328), .Y(n2402) );
  NAND2X1 U1139 ( .A(n1329), .B(n1330), .Y(n1317) );
  NOR2X1 U1140 ( .A(n1318), .B(n1328), .Y(n2403) );
  NAND2X1 U1141 ( .A(n1329), .B(n1331), .Y(n1318) );
  NOR2X1 U1142 ( .A(n1319), .B(n1328), .Y(n2404) );
  NAND2X1 U1143 ( .A(n1329), .B(n1332), .Y(n1319) );
  NOR2X1 U1144 ( .A(n1320), .B(n1328), .Y(n2405) );
  NAND2X1 U1145 ( .A(n1329), .B(n1333), .Y(n1320) );
  NOR2X1 U1146 ( .A(n228), .B(n229), .Y(n1329) );
  NOR2X1 U1147 ( .A(n1321), .B(n1328), .Y(n2406) );
  NOR2X1 U1148 ( .A(n1304), .B(n1328), .Y(n2407) );
  NAND2X1 U1149 ( .A(n1331), .B(n1334), .Y(n1304) );
  NOR2X1 U1150 ( .A(n1305), .B(n1328), .Y(n2408) );
  NAND2X1 U1151 ( .A(n1332), .B(n1334), .Y(n1305) );
  NOR2X1 U1152 ( .A(n1306), .B(n1328), .Y(n2409) );
  NAND2X1 U1153 ( .A(n1333), .B(n1334), .Y(n1306) );
  NOR2X1 U1154 ( .A(n1307), .B(n1328), .Y(n2410) );
  NAND2X1 U1155 ( .A(n1335), .B(n1330), .Y(n1307) );
  NOR2X1 U1156 ( .A(n1308), .B(n1328), .Y(n2411) );
  NAND2X1 U1157 ( .A(n1335), .B(n1331), .Y(n1308) );
  NOR2X1 U1158 ( .A(n1309), .B(n1328), .Y(n2412) );
  NAND2X1 U1159 ( .A(n1335), .B(n1332), .Y(n1309) );
  NOR2X1 U1160 ( .A(n1310), .B(n1328), .Y(n2413) );
  NAND2X1 U1161 ( .A(n1335), .B(n1333), .Y(n1310) );
  NOR2X1 U1162 ( .A(img_counter[3]), .B(n229), .Y(n1335) );
  NOR2X1 U1163 ( .A(n1311), .B(n1328), .Y(n2414) );
  NOR2X1 U1164 ( .A(n1312), .B(n1328), .Y(n2415) );
  NAND2X1 U1165 ( .A(n1331), .B(n1336), .Y(n1312) );
  NOR2X1 U1166 ( .A(img_counter[0]), .B(n230), .Y(n1331) );
  NOR2X1 U1167 ( .A(n1313), .B(n1328), .Y(n2416) );
  NAND2X1 U1168 ( .A(n1332), .B(n1336), .Y(n1313) );
  NOR2X1 U1169 ( .A(img_counter[1]), .B(n231), .Y(n1332) );
  NOR2X1 U1170 ( .A(n1314), .B(n1328), .Y(n2417) );
  NAND3X1 U1171 ( .A(n1315), .B(n225), .C(n226), .Y(n1328) );
  NOR2BX1 U1172 ( .AN(n1325), .B(img_counter[4]), .Y(n1315) );
  AND3X1 U1173 ( .A(n1337), .B(n224), .C(n1338), .Y(n1325) );
  NAND2X1 U1174 ( .A(n1333), .B(n1336), .Y(n1314) );
  NOR2X1 U1175 ( .A(img_counter[0]), .B(img_counter[1]), .Y(n1333) );
  OAI22XL U1176 ( .A0(n431), .A1(n1339), .B0(n1340), .B1(n1341), .Y(n1281) );
  CLKINVX1 U1177 ( .A(n1342), .Y(n1340) );
  OAI211X1 U1178 ( .A0(n1343), .A1(n1344), .B0(n1345), .C0(n1346), .Y(n1342)
         );
  OAI21XL U1179 ( .A0(n1341), .A1(n1347), .B0(n1348), .Y(n1280) );
  MXI2X1 U1180 ( .A(n1349), .B(n1350), .S0(n430), .Y(n1348) );
  NOR2X1 U1181 ( .A(n1341), .B(n1345), .Y(n1350) );
  NAND3BX1 U1182 ( .AN(n1351), .B(n1352), .C(n431), .Y(n1345) );
  OAI21XL U1183 ( .A0(n1353), .A1(n1341), .B0(n1354), .Y(n1279) );
  AO21X1 U1184 ( .A0(n430), .A1(n1355), .B0(n429), .Y(n1354) );
  CLKINVX1 U1185 ( .A(n1349), .Y(n1355) );
  OAI21XL U1186 ( .A0(n431), .A1(n1356), .B0(n1339), .Y(n1349) );
  AOI221XL U1187 ( .A0(n1352), .A1(n1351), .B0(n1357), .B1(n1358), .C0(n1341), 
        .Y(n1339) );
  CLKINVX1 U1188 ( .A(n1344), .Y(n1357) );
  CLKINVX1 U1189 ( .A(n1356), .Y(n1352) );
  OAI21XL U1190 ( .A0(n1359), .A1(n1360), .B0(n1284), .Y(n1341) );
  CLKINVX1 U1191 ( .A(n1361), .Y(n1353) );
  OAI221XL U1192 ( .A0(n1362), .A1(n1363), .B0(n224), .B1(n1364), .C0(n1365), 
        .Y(n1278) );
  NAND2X1 U1193 ( .A(N1167), .B(n1366), .Y(n1365) );
  NAND2X1 U1194 ( .A(n1367), .B(n1368), .Y(n1277) );
  MXI2X1 U1195 ( .A(n1283), .B(cmd[2]), .S0(n1369), .Y(n1367) );
  OAI2BB2XL U1196 ( .B0(n231), .B1(n1364), .A0N(N1160), .A1N(n1366), .Y(n1276)
         );
  OAI2BB2XL U1197 ( .B0(n230), .B1(n1364), .A0N(N1161), .A1N(n1366), .Y(n1275)
         );
  OAI2BB2XL U1198 ( .B0(n229), .B1(n1364), .A0N(N1162), .A1N(n1366), .Y(n1274)
         );
  OAI2BB2XL U1199 ( .B0(n228), .B1(n1364), .A0N(N1163), .A1N(n1366), .Y(n1273)
         );
  OAI221XL U1200 ( .A0(n1343), .A1(n1363), .B0(n227), .B1(n1364), .C0(n1370), 
        .Y(n1272) );
  NAND2X1 U1201 ( .A(N1164), .B(n1366), .Y(n1370) );
  OAI21XL U1202 ( .A0(n226), .A1(n1364), .B0(n1371), .Y(n1271) );
  AOI2BB2X1 U1203 ( .B0(N1165), .B1(n1366), .A0N(n1363), .A1N(n1347), .Y(n1371) );
  OAI221XL U1204 ( .A0(n1363), .A1(n1372), .B0(n225), .B1(n1364), .C0(n1373), 
        .Y(n1270) );
  NAND2X1 U1205 ( .A(N1166), .B(n1366), .Y(n1373) );
  CLKINVX1 U1206 ( .A(n1374), .Y(n1366) );
  AOI32X1 U1207 ( .A0(n1337), .A1(n1284), .A2(n1375), .B0(n1311), .B1(n1376), 
        .Y(n1374) );
  CLKINVX1 U1208 ( .A(n1377), .Y(n1337) );
  NAND3X1 U1209 ( .A(n1378), .B(n1284), .C(n1377), .Y(n1364) );
  NAND2BX1 U1210 ( .AN(n1311), .B(n1376), .Y(n1363) );
  NAND2X1 U1211 ( .A(n1379), .B(n1368), .Y(n1269) );
  MXI2X1 U1212 ( .A(n1285), .B(cmd[0]), .S0(n1369), .Y(n1379) );
  NAND2X1 U1213 ( .A(n1380), .B(n1368), .Y(n1268) );
  NAND2X1 U1214 ( .A(n1369), .B(n1284), .Y(n1368) );
  MXI2X1 U1215 ( .A(n1282), .B(cmd[1]), .S0(n1369), .Y(n1380) );
  NAND2X1 U1216 ( .A(n1302), .B(n1381), .Y(n1369) );
  OAI31XL U1217 ( .A0(n1382), .A1(n1360), .A2(n1383), .B0(n1284), .Y(n1381) );
  NAND3X1 U1218 ( .A(n1346), .B(n1375), .C(n217), .Y(n1382) );
  OAI21XL U1219 ( .A0(n205), .A1(n2303), .B0(n1384), .Y(n1267) );
  CLKINVX1 U1220 ( .A(n1376), .Y(n1384) );
  OAI21XL U1221 ( .A0(n2302), .A1(n1385), .B0(n1302), .Y(n1266) );
  NAND2X1 U1222 ( .A(n205), .B(cmd_valid), .Y(n1302) );
  NOR2X1 U1223 ( .A(n1301), .B(n205), .Y(n1385) );
  NAND4X1 U1224 ( .A(n225), .B(n224), .C(n1386), .D(n1387), .Y(n1301) );
  NOR2X1 U1225 ( .A(n227), .B(n226), .Y(n1386) );
  OAI22XL U1226 ( .A0(n1388), .A1(n1286), .B0(n1389), .B1(n1390), .Y(n1265) );
  AOI2BB1X1 U1227 ( .A0N(n1391), .A1N(n1343), .B0(n1392), .Y(n1390) );
  OAI22XL U1228 ( .A0(n426), .A1(n1393), .B0(n1394), .B1(n1389), .Y(n1264) );
  AOI211X1 U1229 ( .A0(n426), .A1(n1392), .B0(n2418), .C0(n1395), .Y(n1394) );
  CLKINVX1 U1230 ( .A(n1347), .Y(n1395) );
  OAI21XL U1231 ( .A0(n1343), .A1(n1396), .B0(n1397), .Y(n1347) );
  OAI22XL U1232 ( .A0(n425), .A1(n1398), .B0(n1399), .B1(n1389), .Y(n1263) );
  AOI31X1 U1233 ( .A0(n426), .A1(n1392), .A2(n425), .B0(n1361), .Y(n1399) );
  NAND2X1 U1234 ( .A(n1372), .B(n1346), .Y(n1361) );
  XOR2X1 U1235 ( .A(n1400), .B(n1397), .Y(n1372) );
  NOR3X1 U1236 ( .A(n1351), .B(n2304), .C(n1401), .Y(n1392) );
  OAI22XL U1237 ( .A0(n1362), .A1(n1389), .B0(n424), .B1(n1402), .Y(n1262) );
  OA21XL U1238 ( .A0(n425), .A1(n1401), .B0(n1398), .Y(n1402) );
  OA21XL U1239 ( .A0(n426), .A1(n1401), .B0(n1393), .Y(n1398) );
  OA21XL U1240 ( .A0(n1286), .A1(n1401), .B0(n1388), .Y(n1393) );
  AOI221XL U1241 ( .A0(n1403), .A1(n1358), .B0(n1351), .B1(n1404), .C0(n1389), 
        .Y(n1388) );
  CLKINVX1 U1242 ( .A(n1401), .Y(n1404) );
  NOR3BXL U1243 ( .AN(n1405), .B(n1406), .C(n1407), .Y(n1351) );
  CLKINVX1 U1244 ( .A(n1408), .Y(n1358) );
  OAI21XL U1245 ( .A0(n1359), .A1(n1383), .B0(n1284), .Y(n1389) );
  CLKINVX1 U1246 ( .A(n1409), .Y(n1359) );
  XNOR2X1 U1247 ( .A(n1410), .B(n1411), .Y(n1362) );
  NOR2BX1 U1248 ( .AN(n1400), .B(n1397), .Y(n1411) );
  NAND2X1 U1249 ( .A(n1396), .B(n1343), .Y(n1397) );
  OAI222XL U1250 ( .A0(n1286), .A1(n1391), .B0(n431), .B1(n1344), .C0(n227), 
        .C1(n1412), .Y(n1343) );
  OAI222XL U1251 ( .A0(n426), .A1(n1391), .B0(n430), .B1(n1344), .C0(n226), 
        .C1(n1412), .Y(n1396) );
  OAI222XL U1252 ( .A0(n425), .A1(n1391), .B0(n429), .B1(n1344), .C0(n225), 
        .C1(n1412), .Y(n1400) );
  OAI22XL U1253 ( .A0(n224), .A1(n1412), .B0(n424), .B1(n1391), .Y(n1410) );
  NAND2X1 U1254 ( .A(n1403), .B(n1408), .Y(n1391) );
  OAI21XL U1255 ( .A0(n1406), .A1(n1413), .B0(n1414), .Y(n1408) );
  OAI21XL U1256 ( .A0(n1415), .A1(n1405), .B0(n1416), .Y(n1414) );
  OAI21XL U1257 ( .A0(n1407), .A1(n1417), .B0(n1344), .Y(n1416) );
  NAND2X1 U1258 ( .A(n1417), .B(n1418), .Y(n1405) );
  OAI22XL U1259 ( .A0(n1419), .A1(n1286), .B0(n431), .B1(n1420), .Y(n1418) );
  OAI22XL U1260 ( .A0(n426), .A1(n1419), .B0(n430), .B1(n1420), .Y(n1417) );
  CLKINVX1 U1261 ( .A(n1407), .Y(n1415) );
  OAI22XL U1262 ( .A0(n425), .A1(n1419), .B0(n429), .B1(n1420), .Y(n1407) );
  CLKINVX1 U1263 ( .A(n1360), .Y(n1420) );
  NAND2X1 U1264 ( .A(n1356), .B(n1344), .Y(n1360) );
  NAND3X1 U1265 ( .A(n1283), .B(n1282), .C(n218), .Y(n1344) );
  NAND3X1 U1266 ( .A(n1283), .B(n1285), .C(n217), .Y(n1356) );
  NOR2X1 U1267 ( .A(n1419), .B(n424), .Y(n1406) );
  CLKINVX1 U1268 ( .A(n1383), .Y(n1419) );
  NAND2X1 U1269 ( .A(n1401), .B(n1413), .Y(n1383) );
  NAND3X1 U1270 ( .A(n217), .B(n1283), .C(n218), .Y(n1401) );
  CLKINVX1 U1271 ( .A(n1413), .Y(n1403) );
  NAND3X1 U1272 ( .A(n1282), .B(n1285), .C(n216), .Y(n1413) );
  CLKINVX1 U1273 ( .A(n1387), .Y(n1412) );
  NOR2X1 U1274 ( .A(n1378), .B(n1311), .Y(n1387) );
  NAND2X1 U1275 ( .A(n1330), .B(n1336), .Y(n1311) );
  NOR2X1 U1276 ( .A(img_counter[2]), .B(img_counter[3]), .Y(n1336) );
  CLKMX2X2 U1277 ( .A(dataout[7]), .B(n1421), .S0(n1376), .Y(n1261) );
  NAND2X1 U1278 ( .A(n1422), .B(n1423), .Y(n1421) );
  NOR4X1 U1279 ( .A(n1424), .B(n1425), .C(n1426), .D(n1427), .Y(n1423) );
  NAND4X1 U1280 ( .A(n1428), .B(n1429), .C(n1430), .D(n1431), .Y(n1427) );
  AOI221XL U1281 ( .A0(n1432), .A1(\img_buff[107][7] ), .B0(n1433), .B1(
        \img_buff[102][7] ), .C0(n1434), .Y(n1431) );
  OAI22XL U1282 ( .A0(n2282), .A1(n1435), .B0(n1436), .B1(n408), .Y(n1434) );
  AOI222XL U1283 ( .A0(n2284), .A1(n1437), .B0(n1438), .B1(\img_buff[103][7] ), 
        .C0(n1439), .C1(\img_buff[101][7] ), .Y(n1430) );
  AOI222XL U1284 ( .A0(n1440), .A1(\img_buff[98][7] ), .B0(n2285), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][7] ), .Y(n1429) );
  AOI222XL U1285 ( .A0(n1443), .A1(\img_buff[94][7] ), .B0(n1444), .B1(
        \img_buff[95][7] ), .C0(n1445), .C1(\img_buff[96][7] ), .Y(n1428) );
  NAND4X1 U1286 ( .A(n1446), .B(n1447), .C(n1448), .D(n1449), .Y(n1426) );
  AOI221XL U1287 ( .A0(n2278), .A1(n1450), .B0(n2279), .B1(n1451), .C0(n1452), 
        .Y(n1449) );
  OAI22XL U1288 ( .A0(n2277), .A1(n1453), .B0(n2276), .B1(n1454), .Y(n1452) );
  AOI222XL U1289 ( .A0(n1455), .A1(\img_buff[87][7] ), .B0(n1456), .B1(
        \img_buff[88][7] ), .C0(n1457), .C1(\img_buff[89][7] ), .Y(n1448) );
  AOI221XL U1290 ( .A0(n1458), .A1(\img_buff[84][7] ), .B0(n1459), .B1(
        \img_buff[82][7] ), .C0(n1460), .Y(n1447) );
  OAI22XL U1291 ( .A0(n2281), .A1(n1461), .B0(n2280), .B1(n1462), .Y(n1460) );
  AOI222XL U1292 ( .A0(n2283), .A1(n1463), .B0(n1464), .B1(\img_buff[83][7] ), 
        .C0(n1465), .C1(\img_buff[81][7] ), .Y(n1446) );
  NAND4X1 U1293 ( .A(n1466), .B(n1467), .C(n1468), .D(n1469), .Y(n1425) );
  AOI221XL U1294 ( .A0(n2272), .A1(n1470), .B0(n1471), .B1(\img_buff[79][7] ), 
        .C0(n1472), .Y(n1469) );
  OAI22XL U1295 ( .A0(n2273), .A1(n1473), .B0(n2270), .B1(n1474), .Y(n1472) );
  AOI222XL U1296 ( .A0(n2274), .A1(n1475), .B0(n1476), .B1(\img_buff[76][7] ), 
        .C0(n1477), .C1(\img_buff[74][7] ), .Y(n1468) );
  AOI222XL U1297 ( .A0(n1478), .A1(\img_buff[73][7] ), .B0(n2275), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][7] ), .Y(n1467) );
  AOI222XL U1298 ( .A0(n1481), .A1(\img_buff[67][7] ), .B0(n1482), .B1(
        \img_buff[68][7] ), .C0(n1483), .C1(\img_buff[69][7] ), .Y(n1466) );
  NAND4X1 U1299 ( .A(n1484), .B(n1485), .C(n1486), .D(n1487), .Y(n1424) );
  AOI221XL U1300 ( .A0(n1488), .A1(\img_buff[63][7] ), .B0(n1489), .B1(
        \img_buff[64][7] ), .C0(n1490), .Y(n1487) );
  OAI22XL U1301 ( .A0(n1491), .A1(n328), .B0(n1492), .B1(n336), .Y(n1490) );
  AOI222XL U1302 ( .A0(n1493), .A1(\img_buff[60][7] ), .B0(n1494), .B1(
        \img_buff[61][7] ), .C0(n1495), .C1(\img_buff[62][7] ), .Y(n1486) );
  AOI221XL U1303 ( .A0(n1496), .A1(\img_buff[57][7] ), .B0(n1497), .B1(
        \img_buff[55][7] ), .C0(n1498), .Y(n1485) );
  OAI22XL U1304 ( .A0(n2269), .A1(n1499), .B0(n2268), .B1(n1500), .Y(n1498) );
  AOI222XL U1305 ( .A0(n2271), .A1(n1501), .B0(n1502), .B1(\img_buff[56][7] ), 
        .C0(n1503), .C1(\img_buff[54][7] ), .Y(n1484) );
  NOR4X1 U1306 ( .A(n1504), .B(n1505), .C(n1506), .D(n1507), .Y(n1422) );
  NAND4X1 U1307 ( .A(n1508), .B(n1509), .C(n1510), .D(n1511), .Y(n1507) );
  AOI221XL U1308 ( .A0(n2298), .A1(n1512), .B0(n1513), .B1(\img_buff[50][7] ), 
        .C0(n1514), .Y(n1511) );
  OAI22XL U1309 ( .A0(n2299), .A1(n1515), .B0(n2296), .B1(n1516), .Y(n1514) );
  AOI222XL U1310 ( .A0(n2300), .A1(n1517), .B0(n1518), .B1(\img_buff[49][7] ), 
        .C0(n1519), .C1(\img_buff[47][7] ), .Y(n1510) );
  AOI222XL U1311 ( .A0(n1520), .A1(\img_buff[44][7] ), .B0(n2301), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][7] ), .Y(n1509) );
  AOI222XL U1312 ( .A0(n1523), .A1(\img_buff[40][7] ), .B0(n1524), .B1(
        \img_buff[41][7] ), .C0(n1525), .C1(\img_buff[42][7] ), .Y(n1508) );
  NAND4X1 U1313 ( .A(n1526), .B(n1527), .C(n1528), .D(n1529), .Y(n1506) );
  AOI221XL U1314 ( .A0(n1530), .A1(\img_buff[38][7] ), .B0(n1531), .B1(
        \img_buff[39][7] ), .C0(n1532), .Y(n1529) );
  OAI22XL U1315 ( .A0(n1533), .A1(n280), .B0(n1534), .B1(n288), .Y(n1532) );
  AOI222XL U1316 ( .A0(n1535), .A1(\img_buff[33][7] ), .B0(n1536), .B1(
        \img_buff[34][7] ), .C0(n1537), .C1(\img_buff[35][7] ), .Y(n1528) );
  AOI221XL U1317 ( .A0(n1538), .A1(\img_buff[30][7] ), .B0(n1539), .B1(
        \img_buff[28][7] ), .C0(n1540), .Y(n1527) );
  OAI22XL U1318 ( .A0(n2295), .A1(n1541), .B0(n2294), .B1(n1542), .Y(n1540) );
  AOI222XL U1319 ( .A0(n2297), .A1(n1543), .B0(n1544), .B1(\img_buff[29][7] ), 
        .C0(n1545), .C1(\img_buff[27][7] ), .Y(n1526) );
  NAND4X1 U1320 ( .A(n1546), .B(n1547), .C(n1548), .D(n1549), .Y(n1505) );
  AOI221XL U1321 ( .A0(n2290), .A1(n1550), .B0(n1551), .B1(\img_buff[23][7] ), 
        .C0(n1552), .Y(n1549) );
  OAI22XL U1322 ( .A0(n2291), .A1(n1553), .B0(n2288), .B1(n1554), .Y(n1552) );
  AOI222XL U1323 ( .A0(n2292), .A1(n1555), .B0(n1556), .B1(\img_buff[22][7] ), 
        .C0(n1557), .C1(\img_buff[20][7] ), .Y(n1548) );
  AOI222XL U1324 ( .A0(n1558), .A1(\img_buff[17][7] ), .B0(n2293), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][7] ), .Y(n1547) );
  AOI222XL U1325 ( .A0(n1561), .A1(\img_buff[13][7] ), .B0(n1562), .B1(
        \img_buff[14][7] ), .C0(n1563), .C1(\img_buff[15][7] ), .Y(n1546) );
  NAND4X1 U1326 ( .A(n1564), .B(n1565), .C(n1566), .D(n1567), .Y(n1504) );
  AOI221XL U1327 ( .A0(n1568), .A1(\img_buff[11][7] ), .B0(n1569), .B1(
        \img_buff[12][7] ), .C0(n1570), .Y(n1567) );
  OAI22XL U1328 ( .A0(n1571), .A1(n232), .B0(n1572), .B1(n240), .Y(n1570) );
  AOI222XL U1329 ( .A0(n1573), .A1(\img_buff[6][7] ), .B0(n1574), .B1(
        \img_buff[7][7] ), .C0(n1575), .C1(\img_buff[8][7] ), .Y(n1566) );
  AOI221XL U1330 ( .A0(n1576), .A1(\img_buff[4][7] ), .B0(n1577), .B1(
        \img_buff[5][7] ), .C0(n1578), .Y(n1565) );
  OAI22XL U1331 ( .A0(n2287), .A1(n1579), .B0(n2286), .B1(n1580), .Y(n1578) );
  AOI222XL U1332 ( .A0(n2289), .A1(n1581), .B0(n1582), .B1(\img_buff[2][7] ), 
        .C0(n1583), .C1(\img_buff[0][7] ), .Y(n1564) );
  CLKMX2X2 U1333 ( .A(dataout[6]), .B(n1584), .S0(n1376), .Y(n1260) );
  NAND2X1 U1334 ( .A(n1585), .B(n1586), .Y(n1584) );
  NOR4X1 U1335 ( .A(n1587), .B(n1588), .C(n1589), .D(n1590), .Y(n1586) );
  NAND4X1 U1336 ( .A(n1591), .B(n1592), .C(n1593), .D(n1594), .Y(n1590) );
  AOI221XL U1337 ( .A0(n1432), .A1(\img_buff[107][6] ), .B0(n1433), .B1(
        \img_buff[102][6] ), .C0(n1595), .Y(n1594) );
  OAI22XL U1338 ( .A0(n2248), .A1(n1435), .B0(n1436), .B1(n409), .Y(n1595) );
  AOI222XL U1339 ( .A0(n2250), .A1(n1437), .B0(n1438), .B1(\img_buff[103][6] ), 
        .C0(n1439), .C1(\img_buff[101][6] ), .Y(n1593) );
  AOI222XL U1340 ( .A0(n1440), .A1(\img_buff[98][6] ), .B0(n2251), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][6] ), .Y(n1592) );
  AOI222XL U1341 ( .A0(n1443), .A1(\img_buff[94][6] ), .B0(n1444), .B1(
        \img_buff[95][6] ), .C0(n1445), .C1(\img_buff[96][6] ), .Y(n1591) );
  NAND4X1 U1342 ( .A(n1596), .B(n1597), .C(n1598), .D(n1599), .Y(n1589) );
  AOI221XL U1343 ( .A0(n2244), .A1(n1450), .B0(n2245), .B1(n1451), .C0(n1600), 
        .Y(n1599) );
  OAI22XL U1344 ( .A0(n2243), .A1(n1453), .B0(n2242), .B1(n1454), .Y(n1600) );
  AOI222XL U1345 ( .A0(n1455), .A1(\img_buff[87][6] ), .B0(n1456), .B1(
        \img_buff[88][6] ), .C0(n1457), .C1(\img_buff[89][6] ), .Y(n1598) );
  AOI221XL U1346 ( .A0(n1458), .A1(\img_buff[84][6] ), .B0(n1459), .B1(
        \img_buff[82][6] ), .C0(n1601), .Y(n1597) );
  OAI22XL U1347 ( .A0(n2247), .A1(n1461), .B0(n2246), .B1(n1462), .Y(n1601) );
  AOI222XL U1348 ( .A0(n2249), .A1(n1463), .B0(n1464), .B1(\img_buff[83][6] ), 
        .C0(n1465), .C1(\img_buff[81][6] ), .Y(n1596) );
  NAND4X1 U1349 ( .A(n1602), .B(n1603), .C(n1604), .D(n1605), .Y(n1588) );
  AOI221XL U1350 ( .A0(n2238), .A1(n1470), .B0(n1471), .B1(\img_buff[79][6] ), 
        .C0(n1606), .Y(n1605) );
  OAI22XL U1351 ( .A0(n2239), .A1(n1473), .B0(n2236), .B1(n1474), .Y(n1606) );
  AOI222XL U1352 ( .A0(n2240), .A1(n1475), .B0(n1476), .B1(\img_buff[76][6] ), 
        .C0(n1477), .C1(\img_buff[74][6] ), .Y(n1604) );
  AOI222XL U1353 ( .A0(n1478), .A1(\img_buff[73][6] ), .B0(n2241), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][6] ), .Y(n1603) );
  AOI222XL U1354 ( .A0(n1481), .A1(\img_buff[67][6] ), .B0(n1482), .B1(
        \img_buff[68][6] ), .C0(n1483), .C1(\img_buff[69][6] ), .Y(n1602) );
  NAND4X1 U1355 ( .A(n1607), .B(n1608), .C(n1609), .D(n1610), .Y(n1587) );
  AOI221XL U1356 ( .A0(n1488), .A1(\img_buff[63][6] ), .B0(n1489), .B1(
        \img_buff[64][6] ), .C0(n1611), .Y(n1610) );
  OAI22XL U1357 ( .A0(n1491), .A1(n329), .B0(n1492), .B1(n337), .Y(n1611) );
  AOI222XL U1358 ( .A0(n1493), .A1(\img_buff[60][6] ), .B0(n1494), .B1(
        \img_buff[61][6] ), .C0(n1495), .C1(\img_buff[62][6] ), .Y(n1609) );
  AOI221XL U1359 ( .A0(n1496), .A1(\img_buff[57][6] ), .B0(n1497), .B1(
        \img_buff[55][6] ), .C0(n1612), .Y(n1608) );
  OAI22XL U1360 ( .A0(n2235), .A1(n1499), .B0(n2234), .B1(n1500), .Y(n1612) );
  AOI222XL U1361 ( .A0(n2237), .A1(n1501), .B0(n1502), .B1(\img_buff[56][6] ), 
        .C0(n1503), .C1(\img_buff[54][6] ), .Y(n1607) );
  NOR4X1 U1362 ( .A(n1613), .B(n1614), .C(n1615), .D(n1616), .Y(n1585) );
  NAND4X1 U1363 ( .A(n1617), .B(n1618), .C(n1619), .D(n1620), .Y(n1616) );
  AOI221XL U1364 ( .A0(n2264), .A1(n1512), .B0(n1513), .B1(\img_buff[50][6] ), 
        .C0(n1621), .Y(n1620) );
  OAI22XL U1365 ( .A0(n2265), .A1(n1515), .B0(n2262), .B1(n1516), .Y(n1621) );
  AOI222XL U1366 ( .A0(n2266), .A1(n1517), .B0(n1518), .B1(\img_buff[49][6] ), 
        .C0(n1519), .C1(\img_buff[47][6] ), .Y(n1619) );
  AOI222XL U1367 ( .A0(n1520), .A1(\img_buff[44][6] ), .B0(n2267), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][6] ), .Y(n1618) );
  AOI222XL U1368 ( .A0(n1523), .A1(\img_buff[40][6] ), .B0(n1524), .B1(
        \img_buff[41][6] ), .C0(n1525), .C1(\img_buff[42][6] ), .Y(n1617) );
  NAND4X1 U1369 ( .A(n1622), .B(n1623), .C(n1624), .D(n1625), .Y(n1615) );
  AOI221XL U1370 ( .A0(n1530), .A1(\img_buff[38][6] ), .B0(n1531), .B1(
        \img_buff[39][6] ), .C0(n1626), .Y(n1625) );
  OAI22XL U1371 ( .A0(n1533), .A1(n281), .B0(n1534), .B1(n289), .Y(n1626) );
  AOI222XL U1372 ( .A0(n1535), .A1(\img_buff[33][6] ), .B0(n1536), .B1(
        \img_buff[34][6] ), .C0(n1537), .C1(\img_buff[35][6] ), .Y(n1624) );
  AOI221XL U1373 ( .A0(n1538), .A1(\img_buff[30][6] ), .B0(n1539), .B1(
        \img_buff[28][6] ), .C0(n1627), .Y(n1623) );
  OAI22XL U1374 ( .A0(n2261), .A1(n1541), .B0(n2260), .B1(n1542), .Y(n1627) );
  AOI222XL U1375 ( .A0(n2263), .A1(n1543), .B0(n1544), .B1(\img_buff[29][6] ), 
        .C0(n1545), .C1(\img_buff[27][6] ), .Y(n1622) );
  NAND4X1 U1376 ( .A(n1628), .B(n1629), .C(n1630), .D(n1631), .Y(n1614) );
  AOI221XL U1377 ( .A0(n2256), .A1(n1550), .B0(n1551), .B1(\img_buff[23][6] ), 
        .C0(n1632), .Y(n1631) );
  OAI22XL U1378 ( .A0(n2257), .A1(n1553), .B0(n2254), .B1(n1554), .Y(n1632) );
  AOI222XL U1379 ( .A0(n2258), .A1(n1555), .B0(n1556), .B1(\img_buff[22][6] ), 
        .C0(n1557), .C1(\img_buff[20][6] ), .Y(n1630) );
  AOI222XL U1380 ( .A0(n1558), .A1(\img_buff[17][6] ), .B0(n2259), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][6] ), .Y(n1629) );
  AOI222XL U1381 ( .A0(n1561), .A1(\img_buff[13][6] ), .B0(n1562), .B1(
        \img_buff[14][6] ), .C0(n1563), .C1(\img_buff[15][6] ), .Y(n1628) );
  NAND4X1 U1382 ( .A(n1633), .B(n1634), .C(n1635), .D(n1636), .Y(n1613) );
  AOI221XL U1383 ( .A0(n1568), .A1(\img_buff[11][6] ), .B0(n1569), .B1(
        \img_buff[12][6] ), .C0(n1637), .Y(n1636) );
  OAI22XL U1384 ( .A0(n1571), .A1(n233), .B0(n1572), .B1(n241), .Y(n1637) );
  AOI222XL U1385 ( .A0(n1573), .A1(\img_buff[6][6] ), .B0(n1574), .B1(
        \img_buff[7][6] ), .C0(n1575), .C1(\img_buff[8][6] ), .Y(n1635) );
  AOI221XL U1386 ( .A0(n1576), .A1(\img_buff[4][6] ), .B0(n1577), .B1(
        \img_buff[5][6] ), .C0(n1638), .Y(n1634) );
  OAI22XL U1387 ( .A0(n2253), .A1(n1579), .B0(n2252), .B1(n1580), .Y(n1638) );
  AOI222XL U1388 ( .A0(n2255), .A1(n1581), .B0(n1582), .B1(\img_buff[2][6] ), 
        .C0(n1583), .C1(\img_buff[0][6] ), .Y(n1633) );
  CLKMX2X2 U1389 ( .A(dataout[5]), .B(n1639), .S0(n1376), .Y(n1259) );
  NAND2X1 U1390 ( .A(n1640), .B(n1641), .Y(n1639) );
  NOR4X1 U1391 ( .A(n1642), .B(n1643), .C(n1644), .D(n1645), .Y(n1641) );
  NAND4X1 U1392 ( .A(n1646), .B(n1647), .C(n1648), .D(n1649), .Y(n1645) );
  AOI221XL U1393 ( .A0(n1432), .A1(\img_buff[107][5] ), .B0(n1433), .B1(
        \img_buff[102][5] ), .C0(n1650), .Y(n1649) );
  OAI22XL U1394 ( .A0(n2214), .A1(n1435), .B0(n1436), .B1(n410), .Y(n1650) );
  AOI222XL U1395 ( .A0(n2216), .A1(n1437), .B0(n1438), .B1(\img_buff[103][5] ), 
        .C0(n1439), .C1(\img_buff[101][5] ), .Y(n1648) );
  AOI222XL U1396 ( .A0(n1440), .A1(\img_buff[98][5] ), .B0(n2217), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][5] ), .Y(n1647) );
  AOI222XL U1397 ( .A0(n1443), .A1(\img_buff[94][5] ), .B0(n1444), .B1(
        \img_buff[95][5] ), .C0(n1445), .C1(\img_buff[96][5] ), .Y(n1646) );
  NAND4X1 U1398 ( .A(n1651), .B(n1652), .C(n1653), .D(n1654), .Y(n1644) );
  AOI221XL U1399 ( .A0(n2210), .A1(n1450), .B0(n2211), .B1(n1451), .C0(n1655), 
        .Y(n1654) );
  OAI22XL U1400 ( .A0(n2209), .A1(n1453), .B0(n2208), .B1(n1454), .Y(n1655) );
  AOI222XL U1401 ( .A0(n1455), .A1(\img_buff[87][5] ), .B0(n1456), .B1(
        \img_buff[88][5] ), .C0(n1457), .C1(\img_buff[89][5] ), .Y(n1653) );
  AOI221XL U1402 ( .A0(n1458), .A1(\img_buff[84][5] ), .B0(n1459), .B1(
        \img_buff[82][5] ), .C0(n1656), .Y(n1652) );
  OAI22XL U1403 ( .A0(n2213), .A1(n1461), .B0(n2212), .B1(n1462), .Y(n1656) );
  AOI222XL U1404 ( .A0(n2215), .A1(n1463), .B0(n1464), .B1(\img_buff[83][5] ), 
        .C0(n1465), .C1(\img_buff[81][5] ), .Y(n1651) );
  NAND4X1 U1405 ( .A(n1657), .B(n1658), .C(n1659), .D(n1660), .Y(n1643) );
  AOI221XL U1406 ( .A0(n2204), .A1(n1470), .B0(n1471), .B1(\img_buff[79][5] ), 
        .C0(n1661), .Y(n1660) );
  OAI22XL U1407 ( .A0(n2205), .A1(n1473), .B0(n2202), .B1(n1474), .Y(n1661) );
  AOI222XL U1408 ( .A0(n2206), .A1(n1475), .B0(n1476), .B1(\img_buff[76][5] ), 
        .C0(n1477), .C1(\img_buff[74][5] ), .Y(n1659) );
  AOI222XL U1409 ( .A0(n1478), .A1(\img_buff[73][5] ), .B0(n2207), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][5] ), .Y(n1658) );
  AOI222XL U1410 ( .A0(n1481), .A1(\img_buff[67][5] ), .B0(n1482), .B1(
        \img_buff[68][5] ), .C0(n1483), .C1(\img_buff[69][5] ), .Y(n1657) );
  NAND4X1 U1411 ( .A(n1662), .B(n1663), .C(n1664), .D(n1665), .Y(n1642) );
  AOI221XL U1412 ( .A0(n1488), .A1(\img_buff[63][5] ), .B0(n1489), .B1(
        \img_buff[64][5] ), .C0(n1666), .Y(n1665) );
  OAI22XL U1413 ( .A0(n1491), .A1(n330), .B0(n1492), .B1(n338), .Y(n1666) );
  AOI222XL U1414 ( .A0(n1493), .A1(\img_buff[60][5] ), .B0(n1494), .B1(
        \img_buff[61][5] ), .C0(n1495), .C1(\img_buff[62][5] ), .Y(n1664) );
  AOI221XL U1415 ( .A0(n1496), .A1(\img_buff[57][5] ), .B0(n1497), .B1(
        \img_buff[55][5] ), .C0(n1667), .Y(n1663) );
  OAI22XL U1416 ( .A0(n2201), .A1(n1499), .B0(n2200), .B1(n1500), .Y(n1667) );
  AOI222XL U1417 ( .A0(n2203), .A1(n1501), .B0(n1502), .B1(\img_buff[56][5] ), 
        .C0(n1503), .C1(\img_buff[54][5] ), .Y(n1662) );
  NOR4X1 U1418 ( .A(n1668), .B(n1669), .C(n1670), .D(n1671), .Y(n1640) );
  NAND4X1 U1419 ( .A(n1672), .B(n1673), .C(n1674), .D(n1675), .Y(n1671) );
  AOI221XL U1420 ( .A0(n2230), .A1(n1512), .B0(n1513), .B1(\img_buff[50][5] ), 
        .C0(n1676), .Y(n1675) );
  OAI22XL U1421 ( .A0(n2231), .A1(n1515), .B0(n2228), .B1(n1516), .Y(n1676) );
  AOI222XL U1422 ( .A0(n2232), .A1(n1517), .B0(n1518), .B1(\img_buff[49][5] ), 
        .C0(n1519), .C1(\img_buff[47][5] ), .Y(n1674) );
  AOI222XL U1423 ( .A0(n1520), .A1(\img_buff[44][5] ), .B0(n2233), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][5] ), .Y(n1673) );
  AOI222XL U1424 ( .A0(n1523), .A1(\img_buff[40][5] ), .B0(n1524), .B1(
        \img_buff[41][5] ), .C0(n1525), .C1(\img_buff[42][5] ), .Y(n1672) );
  NAND4X1 U1425 ( .A(n1677), .B(n1678), .C(n1679), .D(n1680), .Y(n1670) );
  AOI221XL U1426 ( .A0(n1530), .A1(\img_buff[38][5] ), .B0(n1531), .B1(
        \img_buff[39][5] ), .C0(n1681), .Y(n1680) );
  OAI22XL U1427 ( .A0(n1533), .A1(n282), .B0(n1534), .B1(n290), .Y(n1681) );
  AOI222XL U1428 ( .A0(n1535), .A1(\img_buff[33][5] ), .B0(n1536), .B1(
        \img_buff[34][5] ), .C0(n1537), .C1(\img_buff[35][5] ), .Y(n1679) );
  AOI221XL U1429 ( .A0(n1538), .A1(\img_buff[30][5] ), .B0(n1539), .B1(
        \img_buff[28][5] ), .C0(n1682), .Y(n1678) );
  OAI22XL U1430 ( .A0(n2227), .A1(n1541), .B0(n2226), .B1(n1542), .Y(n1682) );
  AOI222XL U1431 ( .A0(n2229), .A1(n1543), .B0(n1544), .B1(\img_buff[29][5] ), 
        .C0(n1545), .C1(\img_buff[27][5] ), .Y(n1677) );
  NAND4X1 U1432 ( .A(n1683), .B(n1684), .C(n1685), .D(n1686), .Y(n1669) );
  AOI221XL U1433 ( .A0(n2222), .A1(n1550), .B0(n1551), .B1(\img_buff[23][5] ), 
        .C0(n1687), .Y(n1686) );
  OAI22XL U1434 ( .A0(n2223), .A1(n1553), .B0(n2220), .B1(n1554), .Y(n1687) );
  AOI222XL U1435 ( .A0(n2224), .A1(n1555), .B0(n1556), .B1(\img_buff[22][5] ), 
        .C0(n1557), .C1(\img_buff[20][5] ), .Y(n1685) );
  AOI222XL U1436 ( .A0(n1558), .A1(\img_buff[17][5] ), .B0(n2225), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][5] ), .Y(n1684) );
  AOI222XL U1437 ( .A0(n1561), .A1(\img_buff[13][5] ), .B0(n1562), .B1(
        \img_buff[14][5] ), .C0(n1563), .C1(\img_buff[15][5] ), .Y(n1683) );
  NAND4X1 U1438 ( .A(n1688), .B(n1689), .C(n1690), .D(n1691), .Y(n1668) );
  AOI221XL U1439 ( .A0(n1568), .A1(\img_buff[11][5] ), .B0(n1569), .B1(
        \img_buff[12][5] ), .C0(n1692), .Y(n1691) );
  OAI22XL U1440 ( .A0(n1571), .A1(n234), .B0(n1572), .B1(n242), .Y(n1692) );
  AOI222XL U1441 ( .A0(n1573), .A1(\img_buff[6][5] ), .B0(n1574), .B1(
        \img_buff[7][5] ), .C0(n1575), .C1(\img_buff[8][5] ), .Y(n1690) );
  AOI221XL U1442 ( .A0(n1576), .A1(\img_buff[4][5] ), .B0(n1577), .B1(
        \img_buff[5][5] ), .C0(n1693), .Y(n1689) );
  OAI22XL U1443 ( .A0(n2219), .A1(n1579), .B0(n2218), .B1(n1580), .Y(n1693) );
  AOI222XL U1444 ( .A0(n2221), .A1(n1581), .B0(n1582), .B1(\img_buff[2][5] ), 
        .C0(n1583), .C1(\img_buff[0][5] ), .Y(n1688) );
  CLKMX2X2 U1445 ( .A(dataout[4]), .B(n1694), .S0(n1376), .Y(n1258) );
  NAND2X1 U1446 ( .A(n1695), .B(n1696), .Y(n1694) );
  NOR4X1 U1447 ( .A(n1697), .B(n1698), .C(n1699), .D(n1700), .Y(n1696) );
  NAND4X1 U1448 ( .A(n1701), .B(n1702), .C(n1703), .D(n1704), .Y(n1700) );
  AOI221XL U1449 ( .A0(n1432), .A1(\img_buff[107][4] ), .B0(n1433), .B1(
        \img_buff[102][4] ), .C0(n1705), .Y(n1704) );
  OAI22XL U1450 ( .A0(n2180), .A1(n1435), .B0(n1436), .B1(n411), .Y(n1705) );
  AOI222XL U1451 ( .A0(n2182), .A1(n1437), .B0(n1438), .B1(\img_buff[103][4] ), 
        .C0(n1439), .C1(\img_buff[101][4] ), .Y(n1703) );
  AOI222XL U1452 ( .A0(n1440), .A1(\img_buff[98][4] ), .B0(n2183), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][4] ), .Y(n1702) );
  AOI222XL U1453 ( .A0(n1443), .A1(\img_buff[94][4] ), .B0(n1444), .B1(
        \img_buff[95][4] ), .C0(n1445), .C1(\img_buff[96][4] ), .Y(n1701) );
  NAND4X1 U1454 ( .A(n1706), .B(n1707), .C(n1708), .D(n1709), .Y(n1699) );
  AOI221XL U1455 ( .A0(n2176), .A1(n1450), .B0(n2177), .B1(n1451), .C0(n1710), 
        .Y(n1709) );
  OAI22XL U1456 ( .A0(n2175), .A1(n1453), .B0(n2174), .B1(n1454), .Y(n1710) );
  AOI222XL U1457 ( .A0(n1455), .A1(\img_buff[87][4] ), .B0(n1456), .B1(
        \img_buff[88][4] ), .C0(n1457), .C1(\img_buff[89][4] ), .Y(n1708) );
  AOI221XL U1458 ( .A0(n1458), .A1(\img_buff[84][4] ), .B0(n1459), .B1(
        \img_buff[82][4] ), .C0(n1711), .Y(n1707) );
  OAI22XL U1459 ( .A0(n2179), .A1(n1461), .B0(n2178), .B1(n1462), .Y(n1711) );
  AOI222XL U1460 ( .A0(n2181), .A1(n1463), .B0(n1464), .B1(\img_buff[83][4] ), 
        .C0(n1465), .C1(\img_buff[81][4] ), .Y(n1706) );
  NAND4X1 U1461 ( .A(n1712), .B(n1713), .C(n1714), .D(n1715), .Y(n1698) );
  AOI221XL U1462 ( .A0(n2170), .A1(n1470), .B0(n1471), .B1(\img_buff[79][4] ), 
        .C0(n1716), .Y(n1715) );
  OAI22XL U1463 ( .A0(n2171), .A1(n1473), .B0(n2168), .B1(n1474), .Y(n1716) );
  AOI222XL U1464 ( .A0(n2172), .A1(n1475), .B0(n1476), .B1(\img_buff[76][4] ), 
        .C0(n1477), .C1(\img_buff[74][4] ), .Y(n1714) );
  AOI222XL U1465 ( .A0(n1478), .A1(\img_buff[73][4] ), .B0(n2173), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][4] ), .Y(n1713) );
  AOI222XL U1466 ( .A0(n1481), .A1(\img_buff[67][4] ), .B0(n1482), .B1(
        \img_buff[68][4] ), .C0(n1483), .C1(\img_buff[69][4] ), .Y(n1712) );
  NAND4X1 U1467 ( .A(n1717), .B(n1718), .C(n1719), .D(n1720), .Y(n1697) );
  AOI221XL U1468 ( .A0(n1488), .A1(\img_buff[63][4] ), .B0(n1489), .B1(
        \img_buff[64][4] ), .C0(n1721), .Y(n1720) );
  OAI22XL U1469 ( .A0(n1491), .A1(n331), .B0(n1492), .B1(n339), .Y(n1721) );
  AOI222XL U1470 ( .A0(n1493), .A1(\img_buff[60][4] ), .B0(n1494), .B1(
        \img_buff[61][4] ), .C0(n1495), .C1(\img_buff[62][4] ), .Y(n1719) );
  AOI221XL U1471 ( .A0(n1496), .A1(\img_buff[57][4] ), .B0(n1497), .B1(
        \img_buff[55][4] ), .C0(n1722), .Y(n1718) );
  OAI22XL U1472 ( .A0(n2167), .A1(n1499), .B0(n2166), .B1(n1500), .Y(n1722) );
  AOI222XL U1473 ( .A0(n2169), .A1(n1501), .B0(n1502), .B1(\img_buff[56][4] ), 
        .C0(n1503), .C1(\img_buff[54][4] ), .Y(n1717) );
  NOR4X1 U1474 ( .A(n1723), .B(n1724), .C(n1725), .D(n1726), .Y(n1695) );
  NAND4X1 U1475 ( .A(n1727), .B(n1728), .C(n1729), .D(n1730), .Y(n1726) );
  AOI221XL U1476 ( .A0(n2196), .A1(n1512), .B0(n1513), .B1(\img_buff[50][4] ), 
        .C0(n1731), .Y(n1730) );
  OAI22XL U1477 ( .A0(n2197), .A1(n1515), .B0(n2194), .B1(n1516), .Y(n1731) );
  AOI222XL U1478 ( .A0(n2198), .A1(n1517), .B0(n1518), .B1(\img_buff[49][4] ), 
        .C0(n1519), .C1(\img_buff[47][4] ), .Y(n1729) );
  AOI222XL U1479 ( .A0(n1520), .A1(\img_buff[44][4] ), .B0(n2199), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][4] ), .Y(n1728) );
  AOI222XL U1480 ( .A0(n1523), .A1(\img_buff[40][4] ), .B0(n1524), .B1(
        \img_buff[41][4] ), .C0(n1525), .C1(\img_buff[42][4] ), .Y(n1727) );
  NAND4X1 U1481 ( .A(n1732), .B(n1733), .C(n1734), .D(n1735), .Y(n1725) );
  AOI221XL U1482 ( .A0(n1530), .A1(\img_buff[38][4] ), .B0(n1531), .B1(
        \img_buff[39][4] ), .C0(n1736), .Y(n1735) );
  OAI22XL U1483 ( .A0(n1533), .A1(n283), .B0(n1534), .B1(n291), .Y(n1736) );
  AOI222XL U1484 ( .A0(n1535), .A1(\img_buff[33][4] ), .B0(n1536), .B1(
        \img_buff[34][4] ), .C0(n1537), .C1(\img_buff[35][4] ), .Y(n1734) );
  AOI221XL U1485 ( .A0(n1538), .A1(\img_buff[30][4] ), .B0(n1539), .B1(
        \img_buff[28][4] ), .C0(n1737), .Y(n1733) );
  OAI22XL U1486 ( .A0(n2193), .A1(n1541), .B0(n2192), .B1(n1542), .Y(n1737) );
  AOI222XL U1487 ( .A0(n2195), .A1(n1543), .B0(n1544), .B1(\img_buff[29][4] ), 
        .C0(n1545), .C1(\img_buff[27][4] ), .Y(n1732) );
  NAND4X1 U1488 ( .A(n1738), .B(n1739), .C(n1740), .D(n1741), .Y(n1724) );
  AOI221XL U1489 ( .A0(n2188), .A1(n1550), .B0(n1551), .B1(\img_buff[23][4] ), 
        .C0(n1742), .Y(n1741) );
  OAI22XL U1490 ( .A0(n2189), .A1(n1553), .B0(n2186), .B1(n1554), .Y(n1742) );
  AOI222XL U1491 ( .A0(n2190), .A1(n1555), .B0(n1556), .B1(\img_buff[22][4] ), 
        .C0(n1557), .C1(\img_buff[20][4] ), .Y(n1740) );
  AOI222XL U1492 ( .A0(n1558), .A1(\img_buff[17][4] ), .B0(n2191), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][4] ), .Y(n1739) );
  AOI222XL U1493 ( .A0(n1561), .A1(\img_buff[13][4] ), .B0(n1562), .B1(
        \img_buff[14][4] ), .C0(n1563), .C1(\img_buff[15][4] ), .Y(n1738) );
  NAND4X1 U1494 ( .A(n1743), .B(n1744), .C(n1745), .D(n1746), .Y(n1723) );
  AOI221XL U1495 ( .A0(n1568), .A1(\img_buff[11][4] ), .B0(n1569), .B1(
        \img_buff[12][4] ), .C0(n1747), .Y(n1746) );
  OAI22XL U1496 ( .A0(n1571), .A1(n235), .B0(n1572), .B1(n243), .Y(n1747) );
  AOI222XL U1497 ( .A0(n1573), .A1(\img_buff[6][4] ), .B0(n1574), .B1(
        \img_buff[7][4] ), .C0(n1575), .C1(\img_buff[8][4] ), .Y(n1745) );
  AOI221XL U1498 ( .A0(n1576), .A1(\img_buff[4][4] ), .B0(n1577), .B1(
        \img_buff[5][4] ), .C0(n1748), .Y(n1744) );
  OAI22XL U1499 ( .A0(n2185), .A1(n1579), .B0(n2184), .B1(n1580), .Y(n1748) );
  AOI222XL U1500 ( .A0(n2187), .A1(n1581), .B0(n1582), .B1(\img_buff[2][4] ), 
        .C0(n1583), .C1(\img_buff[0][4] ), .Y(n1743) );
  CLKMX2X2 U1501 ( .A(dataout[3]), .B(n1749), .S0(n1376), .Y(n1257) );
  NAND2X1 U1502 ( .A(n1750), .B(n1751), .Y(n1749) );
  NOR4X1 U1503 ( .A(n1752), .B(n1753), .C(n1754), .D(n1755), .Y(n1751) );
  NAND4X1 U1504 ( .A(n1756), .B(n1757), .C(n1758), .D(n1759), .Y(n1755) );
  AOI221XL U1505 ( .A0(n1432), .A1(\img_buff[107][3] ), .B0(n1433), .B1(
        \img_buff[102][3] ), .C0(n1760), .Y(n1759) );
  OAI22XL U1506 ( .A0(n2146), .A1(n1435), .B0(n1436), .B1(n412), .Y(n1760) );
  AOI222XL U1507 ( .A0(n2148), .A1(n1437), .B0(n1438), .B1(\img_buff[103][3] ), 
        .C0(n1439), .C1(\img_buff[101][3] ), .Y(n1758) );
  AOI222XL U1508 ( .A0(n1440), .A1(\img_buff[98][3] ), .B0(n2149), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][3] ), .Y(n1757) );
  AOI222XL U1509 ( .A0(n1443), .A1(\img_buff[94][3] ), .B0(n1444), .B1(
        \img_buff[95][3] ), .C0(n1445), .C1(\img_buff[96][3] ), .Y(n1756) );
  NAND4X1 U1510 ( .A(n1761), .B(n1762), .C(n1763), .D(n1764), .Y(n1754) );
  AOI221XL U1511 ( .A0(n2142), .A1(n1450), .B0(n2143), .B1(n1451), .C0(n1765), 
        .Y(n1764) );
  OAI22XL U1512 ( .A0(n2141), .A1(n1453), .B0(n2140), .B1(n1454), .Y(n1765) );
  AOI222XL U1513 ( .A0(n1455), .A1(\img_buff[87][3] ), .B0(n1456), .B1(
        \img_buff[88][3] ), .C0(n1457), .C1(\img_buff[89][3] ), .Y(n1763) );
  AOI221XL U1514 ( .A0(n1458), .A1(\img_buff[84][3] ), .B0(n1459), .B1(
        \img_buff[82][3] ), .C0(n1766), .Y(n1762) );
  OAI22XL U1515 ( .A0(n2145), .A1(n1461), .B0(n2144), .B1(n1462), .Y(n1766) );
  AOI222XL U1516 ( .A0(n2147), .A1(n1463), .B0(n1464), .B1(\img_buff[83][3] ), 
        .C0(n1465), .C1(\img_buff[81][3] ), .Y(n1761) );
  NAND4X1 U1517 ( .A(n1767), .B(n1768), .C(n1769), .D(n1770), .Y(n1753) );
  AOI221XL U1518 ( .A0(n2136), .A1(n1470), .B0(n1471), .B1(\img_buff[79][3] ), 
        .C0(n1771), .Y(n1770) );
  OAI22XL U1519 ( .A0(n2137), .A1(n1473), .B0(n2134), .B1(n1474), .Y(n1771) );
  AOI222XL U1520 ( .A0(n2138), .A1(n1475), .B0(n1476), .B1(\img_buff[76][3] ), 
        .C0(n1477), .C1(\img_buff[74][3] ), .Y(n1769) );
  AOI222XL U1521 ( .A0(n1478), .A1(\img_buff[73][3] ), .B0(n2139), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][3] ), .Y(n1768) );
  AOI222XL U1522 ( .A0(n1481), .A1(\img_buff[67][3] ), .B0(n1482), .B1(
        \img_buff[68][3] ), .C0(n1483), .C1(\img_buff[69][3] ), .Y(n1767) );
  NAND4X1 U1523 ( .A(n1772), .B(n1773), .C(n1774), .D(n1775), .Y(n1752) );
  AOI221XL U1524 ( .A0(n1488), .A1(\img_buff[63][3] ), .B0(n1489), .B1(
        \img_buff[64][3] ), .C0(n1776), .Y(n1775) );
  OAI22XL U1525 ( .A0(n1491), .A1(n332), .B0(n1492), .B1(n340), .Y(n1776) );
  AOI222XL U1526 ( .A0(n1493), .A1(\img_buff[60][3] ), .B0(n1494), .B1(
        \img_buff[61][3] ), .C0(n1495), .C1(\img_buff[62][3] ), .Y(n1774) );
  AOI221XL U1527 ( .A0(n1496), .A1(\img_buff[57][3] ), .B0(n1497), .B1(
        \img_buff[55][3] ), .C0(n1777), .Y(n1773) );
  OAI22XL U1528 ( .A0(n2133), .A1(n1499), .B0(n2132), .B1(n1500), .Y(n1777) );
  AOI222XL U1529 ( .A0(n2135), .A1(n1501), .B0(n1502), .B1(\img_buff[56][3] ), 
        .C0(n1503), .C1(\img_buff[54][3] ), .Y(n1772) );
  NOR4X1 U1530 ( .A(n1778), .B(n1779), .C(n1780), .D(n1781), .Y(n1750) );
  NAND4X1 U1531 ( .A(n1782), .B(n1783), .C(n1784), .D(n1785), .Y(n1781) );
  AOI221XL U1532 ( .A0(n2162), .A1(n1512), .B0(n1513), .B1(\img_buff[50][3] ), 
        .C0(n1786), .Y(n1785) );
  OAI22XL U1533 ( .A0(n2163), .A1(n1515), .B0(n2160), .B1(n1516), .Y(n1786) );
  AOI222XL U1534 ( .A0(n2164), .A1(n1517), .B0(n1518), .B1(\img_buff[49][3] ), 
        .C0(n1519), .C1(\img_buff[47][3] ), .Y(n1784) );
  AOI222XL U1535 ( .A0(n1520), .A1(\img_buff[44][3] ), .B0(n2165), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][3] ), .Y(n1783) );
  AOI222XL U1536 ( .A0(n1523), .A1(\img_buff[40][3] ), .B0(n1524), .B1(
        \img_buff[41][3] ), .C0(n1525), .C1(\img_buff[42][3] ), .Y(n1782) );
  NAND4X1 U1537 ( .A(n1787), .B(n1788), .C(n1789), .D(n1790), .Y(n1780) );
  AOI221XL U1538 ( .A0(n1530), .A1(\img_buff[38][3] ), .B0(n1531), .B1(
        \img_buff[39][3] ), .C0(n1791), .Y(n1790) );
  OAI22XL U1539 ( .A0(n1533), .A1(n284), .B0(n1534), .B1(n292), .Y(n1791) );
  AOI222XL U1540 ( .A0(n1535), .A1(\img_buff[33][3] ), .B0(n1536), .B1(
        \img_buff[34][3] ), .C0(n1537), .C1(\img_buff[35][3] ), .Y(n1789) );
  AOI221XL U1541 ( .A0(n1538), .A1(\img_buff[30][3] ), .B0(n1539), .B1(
        \img_buff[28][3] ), .C0(n1792), .Y(n1788) );
  OAI22XL U1542 ( .A0(n2159), .A1(n1541), .B0(n2158), .B1(n1542), .Y(n1792) );
  AOI222XL U1543 ( .A0(n2161), .A1(n1543), .B0(n1544), .B1(\img_buff[29][3] ), 
        .C0(n1545), .C1(\img_buff[27][3] ), .Y(n1787) );
  NAND4X1 U1544 ( .A(n1793), .B(n1794), .C(n1795), .D(n1796), .Y(n1779) );
  AOI221XL U1545 ( .A0(n2154), .A1(n1550), .B0(n1551), .B1(\img_buff[23][3] ), 
        .C0(n1797), .Y(n1796) );
  OAI22XL U1546 ( .A0(n2155), .A1(n1553), .B0(n2152), .B1(n1554), .Y(n1797) );
  AOI222XL U1547 ( .A0(n2156), .A1(n1555), .B0(n1556), .B1(\img_buff[22][3] ), 
        .C0(n1557), .C1(\img_buff[20][3] ), .Y(n1795) );
  AOI222XL U1548 ( .A0(n1558), .A1(\img_buff[17][3] ), .B0(n2157), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][3] ), .Y(n1794) );
  AOI222XL U1549 ( .A0(n1561), .A1(\img_buff[13][3] ), .B0(n1562), .B1(
        \img_buff[14][3] ), .C0(n1563), .C1(\img_buff[15][3] ), .Y(n1793) );
  NAND4X1 U1550 ( .A(n1798), .B(n1799), .C(n1800), .D(n1801), .Y(n1778) );
  AOI221XL U1551 ( .A0(n1568), .A1(\img_buff[11][3] ), .B0(n1569), .B1(
        \img_buff[12][3] ), .C0(n1802), .Y(n1801) );
  OAI22XL U1552 ( .A0(n1571), .A1(n236), .B0(n1572), .B1(n244), .Y(n1802) );
  AOI222XL U1553 ( .A0(n1573), .A1(\img_buff[6][3] ), .B0(n1574), .B1(
        \img_buff[7][3] ), .C0(n1575), .C1(\img_buff[8][3] ), .Y(n1800) );
  AOI221XL U1554 ( .A0(n1576), .A1(\img_buff[4][3] ), .B0(n1577), .B1(
        \img_buff[5][3] ), .C0(n1803), .Y(n1799) );
  OAI22XL U1555 ( .A0(n2151), .A1(n1579), .B0(n2150), .B1(n1580), .Y(n1803) );
  AOI222XL U1556 ( .A0(n2153), .A1(n1581), .B0(n1582), .B1(\img_buff[2][3] ), 
        .C0(n1583), .C1(\img_buff[0][3] ), .Y(n1798) );
  CLKMX2X2 U1557 ( .A(dataout[2]), .B(n1804), .S0(n1376), .Y(n1256) );
  NAND2X1 U1558 ( .A(n1805), .B(n1806), .Y(n1804) );
  NOR4X1 U1559 ( .A(n1807), .B(n1808), .C(n1809), .D(n1810), .Y(n1806) );
  NAND4X1 U1560 ( .A(n1811), .B(n1812), .C(n1813), .D(n1814), .Y(n1810) );
  AOI221XL U1561 ( .A0(n1432), .A1(\img_buff[107][2] ), .B0(n1433), .B1(
        \img_buff[102][2] ), .C0(n1815), .Y(n1814) );
  OAI22XL U1562 ( .A0(n2112), .A1(n1435), .B0(n1436), .B1(n413), .Y(n1815) );
  AOI222XL U1563 ( .A0(n2114), .A1(n1437), .B0(n1438), .B1(\img_buff[103][2] ), 
        .C0(n1439), .C1(\img_buff[101][2] ), .Y(n1813) );
  AOI222XL U1564 ( .A0(n1440), .A1(\img_buff[98][2] ), .B0(n2115), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][2] ), .Y(n1812) );
  AOI222XL U1565 ( .A0(n1443), .A1(\img_buff[94][2] ), .B0(n1444), .B1(
        \img_buff[95][2] ), .C0(n1445), .C1(\img_buff[96][2] ), .Y(n1811) );
  NAND4X1 U1566 ( .A(n1816), .B(n1817), .C(n1818), .D(n1819), .Y(n1809) );
  AOI221XL U1567 ( .A0(n2108), .A1(n1450), .B0(n2109), .B1(n1451), .C0(n1820), 
        .Y(n1819) );
  OAI22XL U1568 ( .A0(n2107), .A1(n1453), .B0(n2106), .B1(n1454), .Y(n1820) );
  AOI222XL U1569 ( .A0(n1455), .A1(\img_buff[87][2] ), .B0(n1456), .B1(
        \img_buff[88][2] ), .C0(n1457), .C1(\img_buff[89][2] ), .Y(n1818) );
  AOI221XL U1570 ( .A0(n1458), .A1(\img_buff[84][2] ), .B0(n1459), .B1(
        \img_buff[82][2] ), .C0(n1821), .Y(n1817) );
  OAI22XL U1571 ( .A0(n2111), .A1(n1461), .B0(n2110), .B1(n1462), .Y(n1821) );
  AOI222XL U1572 ( .A0(n2113), .A1(n1463), .B0(n1464), .B1(\img_buff[83][2] ), 
        .C0(n1465), .C1(\img_buff[81][2] ), .Y(n1816) );
  NAND4X1 U1573 ( .A(n1822), .B(n1823), .C(n1824), .D(n1825), .Y(n1808) );
  AOI221XL U1574 ( .A0(n2102), .A1(n1470), .B0(n1471), .B1(\img_buff[79][2] ), 
        .C0(n1826), .Y(n1825) );
  OAI22XL U1575 ( .A0(n2103), .A1(n1473), .B0(n2100), .B1(n1474), .Y(n1826) );
  AOI222XL U1576 ( .A0(n2104), .A1(n1475), .B0(n1476), .B1(\img_buff[76][2] ), 
        .C0(n1477), .C1(\img_buff[74][2] ), .Y(n1824) );
  AOI222XL U1577 ( .A0(n1478), .A1(\img_buff[73][2] ), .B0(n2105), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][2] ), .Y(n1823) );
  AOI222XL U1578 ( .A0(n1481), .A1(\img_buff[67][2] ), .B0(n1482), .B1(
        \img_buff[68][2] ), .C0(n1483), .C1(\img_buff[69][2] ), .Y(n1822) );
  NAND4X1 U1579 ( .A(n1827), .B(n1828), .C(n1829), .D(n1830), .Y(n1807) );
  AOI221XL U1580 ( .A0(n1488), .A1(\img_buff[63][2] ), .B0(n1489), .B1(
        \img_buff[64][2] ), .C0(n1831), .Y(n1830) );
  OAI22XL U1581 ( .A0(n1491), .A1(n333), .B0(n1492), .B1(n341), .Y(n1831) );
  AOI222XL U1582 ( .A0(n1493), .A1(\img_buff[60][2] ), .B0(n1494), .B1(
        \img_buff[61][2] ), .C0(n1495), .C1(\img_buff[62][2] ), .Y(n1829) );
  AOI221XL U1583 ( .A0(n1496), .A1(\img_buff[57][2] ), .B0(n1497), .B1(
        \img_buff[55][2] ), .C0(n1832), .Y(n1828) );
  OAI22XL U1584 ( .A0(n2099), .A1(n1499), .B0(n2098), .B1(n1500), .Y(n1832) );
  AOI222XL U1585 ( .A0(n2101), .A1(n1501), .B0(n1502), .B1(\img_buff[56][2] ), 
        .C0(n1503), .C1(\img_buff[54][2] ), .Y(n1827) );
  NOR4X1 U1586 ( .A(n1833), .B(n1834), .C(n1835), .D(n1836), .Y(n1805) );
  NAND4X1 U1587 ( .A(n1837), .B(n1838), .C(n1839), .D(n1840), .Y(n1836) );
  AOI221XL U1588 ( .A0(n2128), .A1(n1512), .B0(n1513), .B1(\img_buff[50][2] ), 
        .C0(n1841), .Y(n1840) );
  OAI22XL U1589 ( .A0(n2129), .A1(n1515), .B0(n2126), .B1(n1516), .Y(n1841) );
  AOI222XL U1590 ( .A0(n2130), .A1(n1517), .B0(n1518), .B1(\img_buff[49][2] ), 
        .C0(n1519), .C1(\img_buff[47][2] ), .Y(n1839) );
  AOI222XL U1591 ( .A0(n1520), .A1(\img_buff[44][2] ), .B0(n2131), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][2] ), .Y(n1838) );
  AOI222XL U1592 ( .A0(n1523), .A1(\img_buff[40][2] ), .B0(n1524), .B1(
        \img_buff[41][2] ), .C0(n1525), .C1(\img_buff[42][2] ), .Y(n1837) );
  NAND4X1 U1593 ( .A(n1842), .B(n1843), .C(n1844), .D(n1845), .Y(n1835) );
  AOI221XL U1594 ( .A0(n1530), .A1(\img_buff[38][2] ), .B0(n1531), .B1(
        \img_buff[39][2] ), .C0(n1846), .Y(n1845) );
  OAI22XL U1595 ( .A0(n1533), .A1(n285), .B0(n1534), .B1(n293), .Y(n1846) );
  AOI222XL U1596 ( .A0(n1535), .A1(\img_buff[33][2] ), .B0(n1536), .B1(
        \img_buff[34][2] ), .C0(n1537), .C1(\img_buff[35][2] ), .Y(n1844) );
  AOI221XL U1597 ( .A0(n1538), .A1(\img_buff[30][2] ), .B0(n1539), .B1(
        \img_buff[28][2] ), .C0(n1847), .Y(n1843) );
  OAI22XL U1598 ( .A0(n2125), .A1(n1541), .B0(n2124), .B1(n1542), .Y(n1847) );
  AOI222XL U1599 ( .A0(n2127), .A1(n1543), .B0(n1544), .B1(\img_buff[29][2] ), 
        .C0(n1545), .C1(\img_buff[27][2] ), .Y(n1842) );
  NAND4X1 U1600 ( .A(n1848), .B(n1849), .C(n1850), .D(n1851), .Y(n1834) );
  AOI221XL U1601 ( .A0(n2120), .A1(n1550), .B0(n1551), .B1(\img_buff[23][2] ), 
        .C0(n1852), .Y(n1851) );
  OAI22XL U1602 ( .A0(n2121), .A1(n1553), .B0(n2118), .B1(n1554), .Y(n1852) );
  AOI222XL U1603 ( .A0(n2122), .A1(n1555), .B0(n1556), .B1(\img_buff[22][2] ), 
        .C0(n1557), .C1(\img_buff[20][2] ), .Y(n1850) );
  AOI222XL U1604 ( .A0(n1558), .A1(\img_buff[17][2] ), .B0(n2123), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][2] ), .Y(n1849) );
  AOI222XL U1605 ( .A0(n1561), .A1(\img_buff[13][2] ), .B0(n1562), .B1(
        \img_buff[14][2] ), .C0(n1563), .C1(\img_buff[15][2] ), .Y(n1848) );
  NAND4X1 U1606 ( .A(n1853), .B(n1854), .C(n1855), .D(n1856), .Y(n1833) );
  AOI221XL U1607 ( .A0(n1568), .A1(\img_buff[11][2] ), .B0(n1569), .B1(
        \img_buff[12][2] ), .C0(n1857), .Y(n1856) );
  OAI22XL U1608 ( .A0(n1571), .A1(n237), .B0(n1572), .B1(n245), .Y(n1857) );
  AOI222XL U1609 ( .A0(n1573), .A1(\img_buff[6][2] ), .B0(n1574), .B1(
        \img_buff[7][2] ), .C0(n1575), .C1(\img_buff[8][2] ), .Y(n1855) );
  AOI221XL U1610 ( .A0(n1576), .A1(\img_buff[4][2] ), .B0(n1577), .B1(
        \img_buff[5][2] ), .C0(n1858), .Y(n1854) );
  OAI22XL U1611 ( .A0(n2117), .A1(n1579), .B0(n2116), .B1(n1580), .Y(n1858) );
  AOI222XL U1612 ( .A0(n2119), .A1(n1581), .B0(n1582), .B1(\img_buff[2][2] ), 
        .C0(n1583), .C1(\img_buff[0][2] ), .Y(n1853) );
  CLKMX2X2 U1613 ( .A(dataout[1]), .B(n1859), .S0(n1376), .Y(n1255) );
  NAND2X1 U1614 ( .A(n1860), .B(n1861), .Y(n1859) );
  NOR4X1 U1615 ( .A(n1862), .B(n1863), .C(n1864), .D(n1865), .Y(n1861) );
  NAND4X1 U1616 ( .A(n1866), .B(n1867), .C(n1868), .D(n1869), .Y(n1865) );
  AOI221XL U1617 ( .A0(n1432), .A1(\img_buff[107][1] ), .B0(n1433), .B1(
        \img_buff[102][1] ), .C0(n1870), .Y(n1869) );
  OAI22XL U1618 ( .A0(n2078), .A1(n1435), .B0(n1436), .B1(n414), .Y(n1870) );
  AOI222XL U1619 ( .A0(n2080), .A1(n1437), .B0(n1438), .B1(\img_buff[103][1] ), 
        .C0(n1439), .C1(\img_buff[101][1] ), .Y(n1868) );
  AOI222XL U1620 ( .A0(n1440), .A1(\img_buff[98][1] ), .B0(n2081), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][1] ), .Y(n1867) );
  AOI222XL U1621 ( .A0(n1443), .A1(\img_buff[94][1] ), .B0(n1444), .B1(
        \img_buff[95][1] ), .C0(n1445), .C1(\img_buff[96][1] ), .Y(n1866) );
  NAND4X1 U1622 ( .A(n1871), .B(n1872), .C(n1873), .D(n1874), .Y(n1864) );
  AOI221XL U1623 ( .A0(n2074), .A1(n1450), .B0(n2075), .B1(n1451), .C0(n1875), 
        .Y(n1874) );
  OAI22XL U1624 ( .A0(n2073), .A1(n1453), .B0(n2072), .B1(n1454), .Y(n1875) );
  AOI222XL U1625 ( .A0(n1455), .A1(\img_buff[87][1] ), .B0(n1456), .B1(
        \img_buff[88][1] ), .C0(n1457), .C1(\img_buff[89][1] ), .Y(n1873) );
  AOI221XL U1626 ( .A0(n1458), .A1(\img_buff[84][1] ), .B0(n1459), .B1(
        \img_buff[82][1] ), .C0(n1876), .Y(n1872) );
  OAI22XL U1627 ( .A0(n2077), .A1(n1461), .B0(n2076), .B1(n1462), .Y(n1876) );
  AOI222XL U1628 ( .A0(n2079), .A1(n1463), .B0(n1464), .B1(\img_buff[83][1] ), 
        .C0(n1465), .C1(\img_buff[81][1] ), .Y(n1871) );
  NAND4X1 U1629 ( .A(n1877), .B(n1878), .C(n1879), .D(n1880), .Y(n1863) );
  AOI221XL U1630 ( .A0(n2068), .A1(n1470), .B0(n1471), .B1(\img_buff[79][1] ), 
        .C0(n1881), .Y(n1880) );
  OAI22XL U1631 ( .A0(n2069), .A1(n1473), .B0(n2066), .B1(n1474), .Y(n1881) );
  AOI222XL U1632 ( .A0(n2070), .A1(n1475), .B0(n1476), .B1(\img_buff[76][1] ), 
        .C0(n1477), .C1(\img_buff[74][1] ), .Y(n1879) );
  AOI222XL U1633 ( .A0(n1478), .A1(\img_buff[73][1] ), .B0(n2071), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][1] ), .Y(n1878) );
  AOI222XL U1634 ( .A0(n1481), .A1(\img_buff[67][1] ), .B0(n1482), .B1(
        \img_buff[68][1] ), .C0(n1483), .C1(\img_buff[69][1] ), .Y(n1877) );
  NAND4X1 U1635 ( .A(n1882), .B(n1883), .C(n1884), .D(n1885), .Y(n1862) );
  AOI221XL U1636 ( .A0(n1488), .A1(\img_buff[63][1] ), .B0(n1489), .B1(
        \img_buff[64][1] ), .C0(n1886), .Y(n1885) );
  OAI22XL U1637 ( .A0(n1491), .A1(n334), .B0(n1492), .B1(n342), .Y(n1886) );
  AOI222XL U1638 ( .A0(n1493), .A1(\img_buff[60][1] ), .B0(n1494), .B1(
        \img_buff[61][1] ), .C0(n1495), .C1(\img_buff[62][1] ), .Y(n1884) );
  AOI221XL U1639 ( .A0(n1496), .A1(\img_buff[57][1] ), .B0(n1497), .B1(
        \img_buff[55][1] ), .C0(n1887), .Y(n1883) );
  OAI22XL U1640 ( .A0(n2065), .A1(n1499), .B0(n2064), .B1(n1500), .Y(n1887) );
  AOI222XL U1641 ( .A0(n2067), .A1(n1501), .B0(n1502), .B1(\img_buff[56][1] ), 
        .C0(n1503), .C1(\img_buff[54][1] ), .Y(n1882) );
  NOR4X1 U1642 ( .A(n1888), .B(n1889), .C(n1890), .D(n1891), .Y(n1860) );
  NAND4X1 U1643 ( .A(n1892), .B(n1893), .C(n1894), .D(n1895), .Y(n1891) );
  AOI221XL U1644 ( .A0(n2094), .A1(n1512), .B0(n1513), .B1(\img_buff[50][1] ), 
        .C0(n1896), .Y(n1895) );
  OAI22XL U1645 ( .A0(n2095), .A1(n1515), .B0(n2092), .B1(n1516), .Y(n1896) );
  AOI222XL U1646 ( .A0(n2096), .A1(n1517), .B0(n1518), .B1(\img_buff[49][1] ), 
        .C0(n1519), .C1(\img_buff[47][1] ), .Y(n1894) );
  AOI222XL U1647 ( .A0(n1520), .A1(\img_buff[44][1] ), .B0(n2097), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][1] ), .Y(n1893) );
  AOI222XL U1648 ( .A0(n1523), .A1(\img_buff[40][1] ), .B0(n1524), .B1(
        \img_buff[41][1] ), .C0(n1525), .C1(\img_buff[42][1] ), .Y(n1892) );
  NAND4X1 U1649 ( .A(n1897), .B(n1898), .C(n1899), .D(n1900), .Y(n1890) );
  AOI221XL U1650 ( .A0(n1530), .A1(\img_buff[38][1] ), .B0(n1531), .B1(
        \img_buff[39][1] ), .C0(n1901), .Y(n1900) );
  OAI22XL U1651 ( .A0(n1533), .A1(n286), .B0(n1534), .B1(n294), .Y(n1901) );
  AOI222XL U1652 ( .A0(n1535), .A1(\img_buff[33][1] ), .B0(n1536), .B1(
        \img_buff[34][1] ), .C0(n1537), .C1(\img_buff[35][1] ), .Y(n1899) );
  AOI221XL U1653 ( .A0(n1538), .A1(\img_buff[30][1] ), .B0(n1539), .B1(
        \img_buff[28][1] ), .C0(n1902), .Y(n1898) );
  OAI22XL U1654 ( .A0(n2091), .A1(n1541), .B0(n2090), .B1(n1542), .Y(n1902) );
  AOI222XL U1655 ( .A0(n2093), .A1(n1543), .B0(n1544), .B1(\img_buff[29][1] ), 
        .C0(n1545), .C1(\img_buff[27][1] ), .Y(n1897) );
  NAND4X1 U1656 ( .A(n1903), .B(n1904), .C(n1905), .D(n1906), .Y(n1889) );
  AOI221XL U1657 ( .A0(n2086), .A1(n1550), .B0(n1551), .B1(\img_buff[23][1] ), 
        .C0(n1907), .Y(n1906) );
  OAI22XL U1658 ( .A0(n2087), .A1(n1553), .B0(n2084), .B1(n1554), .Y(n1907) );
  AOI222XL U1659 ( .A0(n2088), .A1(n1555), .B0(n1556), .B1(\img_buff[22][1] ), 
        .C0(n1557), .C1(\img_buff[20][1] ), .Y(n1905) );
  AOI222XL U1660 ( .A0(n1558), .A1(\img_buff[17][1] ), .B0(n2089), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][1] ), .Y(n1904) );
  AOI222XL U1661 ( .A0(n1561), .A1(\img_buff[13][1] ), .B0(n1562), .B1(
        \img_buff[14][1] ), .C0(n1563), .C1(\img_buff[15][1] ), .Y(n1903) );
  NAND4X1 U1662 ( .A(n1908), .B(n1909), .C(n1910), .D(n1911), .Y(n1888) );
  AOI221XL U1663 ( .A0(n1568), .A1(\img_buff[11][1] ), .B0(n1569), .B1(
        \img_buff[12][1] ), .C0(n1912), .Y(n1911) );
  OAI22XL U1664 ( .A0(n1571), .A1(n238), .B0(n1572), .B1(n246), .Y(n1912) );
  AOI222XL U1665 ( .A0(n1573), .A1(\img_buff[6][1] ), .B0(n1574), .B1(
        \img_buff[7][1] ), .C0(n1575), .C1(\img_buff[8][1] ), .Y(n1910) );
  AOI221XL U1666 ( .A0(n1576), .A1(\img_buff[4][1] ), .B0(n1577), .B1(
        \img_buff[5][1] ), .C0(n1913), .Y(n1909) );
  OAI22XL U1667 ( .A0(n2083), .A1(n1579), .B0(n2082), .B1(n1580), .Y(n1913) );
  AOI222XL U1668 ( .A0(n2085), .A1(n1581), .B0(n1582), .B1(\img_buff[2][1] ), 
        .C0(n1583), .C1(\img_buff[0][1] ), .Y(n1908) );
  CLKMX2X2 U1669 ( .A(dataout[0]), .B(n1914), .S0(n1376), .Y(n1254) );
  NOR2X1 U1670 ( .A(n1378), .B(n205), .Y(n1376) );
  NAND3X1 U1671 ( .A(n1282), .B(n1285), .C(n1283), .Y(n1378) );
  NAND2X1 U1672 ( .A(n1915), .B(n1916), .Y(n1914) );
  NOR4X1 U1673 ( .A(n1917), .B(n1918), .C(n1919), .D(n1920), .Y(n1916) );
  NAND4X1 U1674 ( .A(n1921), .B(n1922), .C(n1923), .D(n1924), .Y(n1920) );
  AOI221XL U1675 ( .A0(n1432), .A1(\img_buff[107][0] ), .B0(n1433), .B1(
        \img_buff[102][0] ), .C0(n1925), .Y(n1924) );
  OAI22XL U1676 ( .A0(n2044), .A1(n1435), .B0(n1436), .B1(n415), .Y(n1925) );
  NAND2X1 U1677 ( .A(n1926), .B(n1927), .Y(n1436) );
  NAND2X1 U1678 ( .A(n1926), .B(n1928), .Y(n1435) );
  AND2X1 U1679 ( .A(n1929), .B(n1928), .Y(n1433) );
  AND2X1 U1680 ( .A(n1926), .B(n1930), .Y(n1432) );
  AOI222XL U1681 ( .A0(n2046), .A1(n1437), .B0(n1438), .B1(\img_buff[103][0] ), 
        .C0(n1439), .C1(\img_buff[101][0] ), .Y(n1923) );
  AND2X1 U1682 ( .A(n1929), .B(n1931), .Y(n1439) );
  AND2X1 U1683 ( .A(n1929), .B(n1930), .Y(n1438) );
  AND2X1 U1684 ( .A(n1929), .B(n1927), .Y(n1437) );
  NOR2BX1 U1685 ( .AN(n1932), .B(n1933), .Y(n1929) );
  AOI222XL U1686 ( .A0(n1440), .A1(\img_buff[98][0] ), .B0(n2047), .B1(n1441), 
        .C0(n1442), .C1(\img_buff[97][0] ), .Y(n1922) );
  AND2X1 U1687 ( .A(n1932), .B(n1934), .Y(n1442) );
  AND2X1 U1688 ( .A(n1932), .B(n1935), .Y(n1441) );
  AND2X1 U1689 ( .A(n1932), .B(n1936), .Y(n1440) );
  AOI222XL U1690 ( .A0(n1443), .A1(\img_buff[94][0] ), .B0(n1444), .B1(
        \img_buff[95][0] ), .C0(n1445), .C1(\img_buff[96][0] ), .Y(n1921) );
  AND2X1 U1691 ( .A(n1932), .B(n1937), .Y(n1445) );
  AND2X1 U1692 ( .A(n1938), .B(n1939), .Y(n1444) );
  AND2X1 U1693 ( .A(n1940), .B(n1939), .Y(n1443) );
  NAND4X1 U1694 ( .A(n1941), .B(n1942), .C(n1943), .D(n1944), .Y(n1919) );
  AOI221XL U1695 ( .A0(n2040), .A1(n1450), .B0(n2041), .B1(n1451), .C0(n1945), 
        .Y(n1944) );
  OAI22XL U1696 ( .A0(n2039), .A1(n1453), .B0(n2038), .B1(n1454), .Y(n1945) );
  NAND2X1 U1697 ( .A(n1946), .B(n1939), .Y(n1454) );
  NAND2X1 U1698 ( .A(n1947), .B(n1939), .Y(n1453) );
  AND2X1 U1699 ( .A(n1940), .B(n1948), .Y(n1451) );
  AND2X1 U1700 ( .A(n1938), .B(n1948), .Y(n1450) );
  AOI222XL U1701 ( .A0(n1455), .A1(\img_buff[87][0] ), .B0(n1456), .B1(
        \img_buff[88][0] ), .C0(n1457), .C1(\img_buff[89][0] ), .Y(n1943) );
  AND2X1 U1702 ( .A(n1947), .B(n1948), .Y(n1457) );
  AND2X1 U1703 ( .A(n1946), .B(n1948), .Y(n1456) );
  AND2X1 U1704 ( .A(n1938), .B(n1949), .Y(n1455) );
  AOI221XL U1705 ( .A0(n1458), .A1(\img_buff[84][0] ), .B0(n1459), .B1(
        \img_buff[82][0] ), .C0(n1950), .Y(n1942) );
  OAI22XL U1706 ( .A0(n2043), .A1(n1461), .B0(n2042), .B1(n1462), .Y(n1950) );
  NAND2X1 U1707 ( .A(n1947), .B(n1949), .Y(n1462) );
  NAND2X1 U1708 ( .A(n1940), .B(n1949), .Y(n1461) );
  AND2X1 U1709 ( .A(n1951), .B(n1940), .Y(n1459) );
  AND2X1 U1710 ( .A(n1946), .B(n1949), .Y(n1458) );
  AOI222XL U1711 ( .A0(n2045), .A1(n1463), .B0(n1464), .B1(\img_buff[83][0] ), 
        .C0(n1465), .C1(\img_buff[81][0] ), .Y(n1941) );
  AND2X1 U1712 ( .A(n1951), .B(n1947), .Y(n1465) );
  AND2X1 U1713 ( .A(n1951), .B(n1938), .Y(n1464) );
  AND2X1 U1714 ( .A(n1926), .B(n1931), .Y(n1463) );
  NOR2BX1 U1715 ( .AN(n1932), .B(n1952), .Y(n1926) );
  NOR2BX1 U1716 ( .AN(out_pos[6]), .B(n1953), .Y(n1932) );
  NAND4X1 U1717 ( .A(n1954), .B(n1955), .C(n1956), .D(n1957), .Y(n1918) );
  AOI221XL U1718 ( .A0(n2034), .A1(n1470), .B0(n1471), .B1(\img_buff[79][0] ), 
        .C0(n1958), .Y(n1957) );
  OAI22XL U1719 ( .A0(n2035), .A1(n1473), .B0(n2032), .B1(n1474), .Y(n1958) );
  NAND2X1 U1720 ( .A(n1951), .B(n1946), .Y(n1474) );
  NAND2X1 U1721 ( .A(n1959), .B(n1930), .Y(n1473) );
  AND2X1 U1722 ( .A(n1938), .B(n1960), .Y(n1471) );
  AND2X1 U1723 ( .A(n1930), .B(out_pos[6]), .Y(n1938) );
  AND2X1 U1724 ( .A(n1947), .B(n1960), .Y(n1470) );
  AND2X1 U1725 ( .A(n1931), .B(out_pos[6]), .Y(n1947) );
  AOI222XL U1726 ( .A0(n2036), .A1(n1475), .B0(n1476), .B1(\img_buff[76][0] ), 
        .C0(n1477), .C1(\img_buff[74][0] ), .Y(n1956) );
  AND2X1 U1727 ( .A(n1959), .B(n1928), .Y(n1477) );
  AND2X1 U1728 ( .A(n1946), .B(n1960), .Y(n1476) );
  AND2X1 U1729 ( .A(n1927), .B(out_pos[6]), .Y(n1946) );
  AND2X1 U1730 ( .A(n1961), .B(n1930), .Y(n1475) );
  AOI222XL U1731 ( .A0(n1478), .A1(\img_buff[73][0] ), .B0(n2037), .B1(n1479), 
        .C0(n1480), .C1(\img_buff[72][0] ), .Y(n1955) );
  AND2X1 U1732 ( .A(n1959), .B(n1927), .Y(n1480) );
  AND2X1 U1733 ( .A(n1961), .B(n1928), .Y(n1479) );
  AND2X1 U1734 ( .A(n1959), .B(n1931), .Y(n1478) );
  AND3X1 U1735 ( .A(out_pos[6]), .B(n1953), .C(n1962), .Y(n1959) );
  AOI222XL U1736 ( .A0(n1481), .A1(\img_buff[67][0] ), .B0(n1482), .B1(
        \img_buff[68][0] ), .C0(n1483), .C1(\img_buff[69][0] ), .Y(n1954) );
  AND2X1 U1737 ( .A(n1961), .B(n1931), .Y(n1483) );
  AND2X1 U1738 ( .A(n1961), .B(n1927), .Y(n1482) );
  AND2X1 U1739 ( .A(n1963), .B(n1964), .Y(n1961) );
  AND2X1 U1740 ( .A(n1935), .B(n1964), .Y(n1481) );
  NAND4X1 U1741 ( .A(n1965), .B(n1966), .C(n1967), .D(n1968), .Y(n1917) );
  AOI221XL U1742 ( .A0(n1488), .A1(\img_buff[63][0] ), .B0(n1489), .B1(
        \img_buff[64][0] ), .C0(n1969), .Y(n1968) );
  OAI22XL U1743 ( .A0(n1491), .A1(n335), .B0(n1492), .B1(n343), .Y(n1969) );
  NAND2X1 U1744 ( .A(n1964), .B(n1936), .Y(n1492) );
  NAND2X1 U1745 ( .A(n1934), .B(n1964), .Y(n1491) );
  AND2X1 U1746 ( .A(n1937), .B(n1964), .Y(n1489) );
  NOR3BXL U1747 ( .AN(out_pos[6]), .B(out_pos[4]), .C(out_pos[5]), .Y(n1964)
         );
  AND2X1 U1748 ( .A(n1970), .B(n1939), .Y(n1488) );
  AOI222XL U1749 ( .A0(n1493), .A1(\img_buff[60][0] ), .B0(n1494), .B1(
        \img_buff[61][0] ), .C0(n1495), .C1(\img_buff[62][0] ), .Y(n1967) );
  AND2X1 U1750 ( .A(n1971), .B(n1939), .Y(n1495) );
  AND2X1 U1751 ( .A(n1972), .B(n1939), .Y(n1494) );
  AND2X1 U1752 ( .A(n1973), .B(n1939), .Y(n1493) );
  AOI221XL U1753 ( .A0(n1496), .A1(\img_buff[57][0] ), .B0(n1497), .B1(
        \img_buff[55][0] ), .C0(n1974), .Y(n1966) );
  OAI22XL U1754 ( .A0(n2031), .A1(n1499), .B0(n2030), .B1(n1500), .Y(n1974) );
  NAND2X1 U1755 ( .A(n1948), .B(n1971), .Y(n1500) );
  NAND2X1 U1756 ( .A(n1948), .B(n1970), .Y(n1499) );
  AND2X1 U1757 ( .A(n1949), .B(n1970), .Y(n1497) );
  AND2X1 U1758 ( .A(n1948), .B(n1972), .Y(n1496) );
  AOI222XL U1759 ( .A0(n2033), .A1(n1501), .B0(n1502), .B1(\img_buff[56][0] ), 
        .C0(n1503), .C1(\img_buff[54][0] ), .Y(n1965) );
  AND2X1 U1760 ( .A(n1949), .B(n1971), .Y(n1503) );
  AND2X1 U1761 ( .A(n1948), .B(n1973), .Y(n1502) );
  AND2X1 U1762 ( .A(n1960), .B(n1940), .Y(n1501) );
  AND2X1 U1763 ( .A(n1928), .B(out_pos[6]), .Y(n1940) );
  NOR4X1 U1764 ( .A(n1975), .B(n1976), .C(n1977), .D(n1978), .Y(n1915) );
  NAND4X1 U1765 ( .A(n1979), .B(n1980), .C(n1981), .D(n1982), .Y(n1978) );
  AOI221XL U1766 ( .A0(n2060), .A1(n1512), .B0(n1513), .B1(\img_buff[50][0] ), 
        .C0(n1983), .Y(n1982) );
  OAI22XL U1767 ( .A0(n2061), .A1(n1515), .B0(n2058), .B1(n1516), .Y(n1983) );
  NAND2X1 U1768 ( .A(n1951), .B(n1970), .Y(n1516) );
  NAND2X1 U1769 ( .A(n1951), .B(n1973), .Y(n1515) );
  AND2X1 U1770 ( .A(n1951), .B(n1971), .Y(n1513) );
  AND2X1 U1771 ( .A(n1949), .B(n1973), .Y(n1512) );
  AOI222XL U1772 ( .A0(n2062), .A1(n1517), .B0(n1518), .B1(\img_buff[49][0] ), 
        .C0(n1519), .C1(\img_buff[47][0] ), .Y(n1981) );
  AND2X1 U1773 ( .A(n1960), .B(n1970), .Y(n1519) );
  NOR2BX1 U1774 ( .AN(n1930), .B(n1953), .Y(n1970) );
  AND2X1 U1775 ( .A(n1951), .B(n1972), .Y(n1518) );
  AND2X1 U1776 ( .A(n1960), .B(n1971), .Y(n1517) );
  NOR2BX1 U1777 ( .AN(n1928), .B(n1953), .Y(n1971) );
  AOI222XL U1778 ( .A0(n1520), .A1(\img_buff[44][0] ), .B0(n2063), .B1(n1521), 
        .C0(n1522), .C1(\img_buff[43][0] ), .Y(n1980) );
  AND2X1 U1779 ( .A(n1984), .B(n1930), .Y(n1522) );
  AND2X1 U1780 ( .A(n1960), .B(n1972), .Y(n1521) );
  AND2X1 U1781 ( .A(n1960), .B(n1973), .Y(n1520) );
  NOR2BX1 U1782 ( .AN(n1927), .B(n1953), .Y(n1973) );
  AOI222XL U1783 ( .A0(n1523), .A1(\img_buff[40][0] ), .B0(n1524), .B1(
        \img_buff[41][0] ), .C0(n1525), .C1(\img_buff[42][0] ), .Y(n1979) );
  AND2X1 U1784 ( .A(n1984), .B(n1928), .Y(n1525) );
  AND2X1 U1785 ( .A(n1984), .B(n1931), .Y(n1524) );
  AND2X1 U1786 ( .A(n1984), .B(n1927), .Y(n1523) );
  NOR3BXL U1787 ( .AN(n1962), .B(n1953), .C(out_pos[6]), .Y(n1984) );
  NAND4X1 U1788 ( .A(n1985), .B(n1986), .C(n1987), .D(n1988), .Y(n1977) );
  AOI221XL U1789 ( .A0(n1530), .A1(\img_buff[38][0] ), .B0(n1531), .B1(
        \img_buff[39][0] ), .C0(n1989), .Y(n1988) );
  OAI22XL U1790 ( .A0(n1533), .A1(n287), .B0(n1534), .B1(n295), .Y(n1989) );
  NAND2X1 U1791 ( .A(n1990), .B(n1931), .Y(n1534) );
  NAND2X1 U1792 ( .A(n1990), .B(n1927), .Y(n1533) );
  AND2X1 U1793 ( .A(n1990), .B(n1930), .Y(n1531) );
  AND2X1 U1794 ( .A(n1990), .B(n1928), .Y(n1530) );
  AND2X1 U1795 ( .A(n1991), .B(n1963), .Y(n1990) );
  AOI222XL U1796 ( .A0(n1535), .A1(\img_buff[33][0] ), .B0(n1536), .B1(
        \img_buff[34][0] ), .C0(n1537), .C1(\img_buff[35][0] ), .Y(n1987) );
  AND2X1 U1797 ( .A(n1991), .B(n1935), .Y(n1537) );
  AND2X1 U1798 ( .A(n1991), .B(n1936), .Y(n1536) );
  AND2X1 U1799 ( .A(n1991), .B(n1934), .Y(n1535) );
  AOI221XL U1800 ( .A0(n1538), .A1(\img_buff[30][0] ), .B0(n1539), .B1(
        \img_buff[28][0] ), .C0(n1992), .Y(n1986) );
  OAI22XL U1801 ( .A0(n2057), .A1(n1541), .B0(n2056), .B1(n1542), .Y(n1992) );
  NAND2X1 U1802 ( .A(n1993), .B(n1939), .Y(n1542) );
  NAND2X1 U1803 ( .A(n1991), .B(n1937), .Y(n1541) );
  NOR3X1 U1804 ( .A(out_pos[4]), .B(out_pos[6]), .C(n1953), .Y(n1991) );
  AND2X1 U1805 ( .A(n1994), .B(n1939), .Y(n1539) );
  AND2X1 U1806 ( .A(n1995), .B(n1939), .Y(n1538) );
  AOI222XL U1807 ( .A0(n2059), .A1(n1543), .B0(n1544), .B1(\img_buff[29][0] ), 
        .C0(n1545), .C1(\img_buff[27][0] ), .Y(n1985) );
  AND2X1 U1808 ( .A(n1993), .B(n1948), .Y(n1545) );
  AND2X1 U1809 ( .A(n1996), .B(n1939), .Y(n1544) );
  NOR3X1 U1810 ( .A(n1952), .B(n1933), .C(n1997), .Y(n1939) );
  AND2X1 U1811 ( .A(n1949), .B(n1972), .Y(n1543) );
  NOR2BX1 U1812 ( .AN(n1931), .B(n1953), .Y(n1972) );
  CLKINVX1 U1813 ( .A(out_pos[5]), .Y(n1953) );
  NAND4X1 U1814 ( .A(n1998), .B(n1999), .C(n2000), .D(n2001), .Y(n1976) );
  AOI221XL U1815 ( .A0(n2052), .A1(n1550), .B0(n1551), .B1(\img_buff[23][0] ), 
        .C0(n2002), .Y(n2001) );
  OAI22XL U1816 ( .A0(n2053), .A1(n1553), .B0(n2050), .B1(n1554), .Y(n2002) );
  NAND2X1 U1817 ( .A(n1994), .B(n1948), .Y(n1554) );
  NAND2X1 U1818 ( .A(n1996), .B(n1949), .Y(n1553) );
  AND2X1 U1819 ( .A(n1993), .B(n1949), .Y(n1551) );
  AND2X1 U1820 ( .A(n1996), .B(n1948), .Y(n1550) );
  AOI222XL U1821 ( .A0(n2054), .A1(n1555), .B0(n1556), .B1(\img_buff[22][0] ), 
        .C0(n1557), .C1(\img_buff[20][0] ), .Y(n2000) );
  AND2X1 U1822 ( .A(n1994), .B(n1949), .Y(n1557) );
  AND2X1 U1823 ( .A(n1995), .B(n1949), .Y(n1556) );
  NOR2BX1 U1824 ( .AN(n1963), .B(n1997), .Y(n1949) );
  AND2X1 U1825 ( .A(n1993), .B(n1951), .Y(n1555) );
  AOI222XL U1826 ( .A0(n1558), .A1(\img_buff[17][0] ), .B0(n2055), .B1(n1559), 
        .C0(n1560), .C1(\img_buff[16][0] ), .Y(n1999) );
  AND2X1 U1827 ( .A(n1994), .B(n1951), .Y(n1560) );
  AND2X1 U1828 ( .A(n1995), .B(n1951), .Y(n1559) );
  AND2X1 U1829 ( .A(n1996), .B(n1951), .Y(n1558) );
  NOR2BX1 U1830 ( .AN(n2003), .B(n1997), .Y(n1951) );
  AOI222XL U1831 ( .A0(n1561), .A1(\img_buff[13][0] ), .B0(n1562), .B1(
        \img_buff[14][0] ), .C0(n1563), .C1(\img_buff[15][0] ), .Y(n1998) );
  AND2X1 U1832 ( .A(n1993), .B(n1960), .Y(n1563) );
  AND2X1 U1833 ( .A(n1995), .B(n1960), .Y(n1562) );
  AND2X1 U1834 ( .A(n1996), .B(n1960), .Y(n1561) );
  NAND4X1 U1835 ( .A(n2004), .B(n2005), .C(n2006), .D(n2007), .Y(n1975) );
  AOI221XL U1836 ( .A0(n1568), .A1(\img_buff[11][0] ), .B0(n1569), .B1(
        \img_buff[12][0] ), .C0(n2008), .Y(n2007) );
  OAI22XL U1837 ( .A0(n1571), .A1(n239), .B0(n1572), .B1(n247), .Y(n2008) );
  NAND2X1 U1838 ( .A(n1995), .B(n1962), .Y(n1572) );
  NAND2X1 U1839 ( .A(n1996), .B(n1962), .Y(n1571) );
  AND2X1 U1840 ( .A(n2009), .B(n1931), .Y(n1996) );
  AND2X1 U1841 ( .A(n1994), .B(n1960), .Y(n1569) );
  NOR3X1 U1842 ( .A(n1933), .B(out_pos[4]), .C(n1952), .Y(n1960) );
  AND2X1 U1843 ( .A(n1993), .B(n1962), .Y(n1568) );
  AND2X1 U1844 ( .A(n2009), .B(n1930), .Y(n1993) );
  AOI222XL U1845 ( .A0(n1573), .A1(\img_buff[6][0] ), .B0(n1574), .B1(
        \img_buff[7][0] ), .C0(n1575), .C1(\img_buff[8][0] ), .Y(n2006) );
  AND2X1 U1846 ( .A(n1994), .B(n1962), .Y(n1575) );
  NOR3X1 U1847 ( .A(out_pos[2]), .B(out_pos[4]), .C(n1952), .Y(n1962) );
  AND2X1 U1848 ( .A(n2009), .B(n1927), .Y(n1994) );
  AND2X1 U1849 ( .A(n2010), .B(n1930), .Y(n1574) );
  AND2X1 U1850 ( .A(n2010), .B(n1928), .Y(n1573) );
  AOI221XL U1851 ( .A0(n1576), .A1(\img_buff[4][0] ), .B0(n1577), .B1(
        \img_buff[5][0] ), .C0(n2011), .Y(n2005) );
  OAI22XL U1852 ( .A0(n2049), .A1(n1579), .B0(n2048), .B1(n1580), .Y(n2011) );
  NAND2X1 U1853 ( .A(n2012), .B(n1935), .Y(n1580) );
  AND2X1 U1854 ( .A(n1930), .B(n2003), .Y(n1935) );
  NOR2BX1 U1855 ( .AN(out_pos[0]), .B(n2013), .Y(n1930) );
  NAND2X1 U1856 ( .A(n2012), .B(n1934), .Y(n1579) );
  AND2X1 U1857 ( .A(n1931), .B(n2003), .Y(n1934) );
  AND2X1 U1858 ( .A(n2010), .B(n1931), .Y(n1577) );
  NOR2BX1 U1859 ( .AN(out_pos[0]), .B(out_pos[1]), .Y(n1931) );
  AND2X1 U1860 ( .A(n2010), .B(n1927), .Y(n1576) );
  AND2X1 U1861 ( .A(n2012), .B(n1963), .Y(n2010) );
  NOR2X1 U1862 ( .A(n1933), .B(out_pos[3]), .Y(n1963) );
  CLKINVX1 U1863 ( .A(out_pos[2]), .Y(n1933) );
  AOI222XL U1864 ( .A0(n2051), .A1(n1581), .B0(n1582), .B1(\img_buff[2][0] ), 
        .C0(n1583), .C1(\img_buff[0][0] ), .Y(n2004) );
  AND2X1 U1865 ( .A(n2012), .B(n1937), .Y(n1583) );
  AND2X1 U1866 ( .A(n1927), .B(n2003), .Y(n1937) );
  NOR2X1 U1867 ( .A(out_pos[0]), .B(out_pos[1]), .Y(n1927) );
  AND2X1 U1868 ( .A(n2012), .B(n1936), .Y(n1582) );
  AND2X1 U1869 ( .A(n1928), .B(n2003), .Y(n1936) );
  NOR2X1 U1870 ( .A(out_pos[2]), .B(out_pos[3]), .Y(n2003) );
  NOR2BX1 U1871 ( .AN(n2009), .B(out_pos[4]), .Y(n2012) );
  AND2X1 U1872 ( .A(n1995), .B(n1948), .Y(n1581) );
  NOR3X1 U1873 ( .A(n1952), .B(out_pos[2]), .C(n1997), .Y(n1948) );
  CLKINVX1 U1874 ( .A(out_pos[4]), .Y(n1997) );
  CLKINVX1 U1875 ( .A(out_pos[3]), .Y(n1952) );
  AND2X1 U1876 ( .A(n2009), .B(n1928), .Y(n1995) );
  NOR2X1 U1877 ( .A(n2013), .B(out_pos[0]), .Y(n1928) );
  CLKINVX1 U1878 ( .A(out_pos[1]), .Y(n2013) );
  NOR2X1 U1879 ( .A(out_pos[5]), .B(out_pos[6]), .Y(n2009) );
  AO21X1 U1880 ( .A0(n1338), .A1(n2014), .B0(n2310), .Y(n1236) );
  NOR3BXL U1881 ( .AN(n1338), .B(n1377), .C(n1375), .Y(n2310) );
  NAND3BX1 U1882 ( .AN(n1321), .B(n2015), .C(n227), .Y(n1375) );
  NOR3BXL U1883 ( .AN(n224), .B(n226), .C(n225), .Y(n2015) );
  NAND2X1 U1884 ( .A(n1334), .B(n1330), .Y(n1321) );
  NOR2X1 U1885 ( .A(n230), .B(n231), .Y(n1330) );
  NOR2X1 U1886 ( .A(img_counter[2]), .B(n228), .Y(n1334) );
  NAND3X1 U1887 ( .A(n217), .B(n216), .C(n218), .Y(n1377) );
  OAI31XL U1888 ( .A0(n1285), .A1(n217), .A2(n1283), .B0(n1409), .Y(n2014) );
  NAND2X1 U1889 ( .A(n2418), .B(n432), .Y(n1409) );
  CLKINVX1 U1890 ( .A(n1346), .Y(n2418) );
  NAND3X1 U1891 ( .A(n216), .B(n1285), .C(n217), .Y(n1346) );
  NOR2X1 U1892 ( .A(n205), .B(reset), .Y(n1338) );
  AND2X1 U1893 ( .A(N973), .B(n432), .Y(\U3/U16/Z_6 ) );
  AND2X1 U1894 ( .A(N972), .B(n432), .Y(\U3/U16/Z_5 ) );
  AND2X1 U1895 ( .A(N971), .B(n432), .Y(\U3/U16/Z_4 ) );
  NOR2X1 U1896 ( .A(n224), .B(n1290), .Y(\U3/U15/Z_6 ) );
  MXI2X1 U1897 ( .A(n2016), .B(n225), .S0(n432), .Y(\U3/U15/Z_5 ) );
  XOR2X1 U1898 ( .A(n2017), .B(n2018), .Y(n2016) );
  NOR2X1 U1899 ( .A(n2019), .B(n2020), .Y(n2018) );
  XOR2X1 U1900 ( .A(n2021), .B(n224), .Y(n2017) );
  OAI22XL U1901 ( .A0(n225), .A1(n2022), .B0(n429), .B1(n2023), .Y(n2021) );
  AND2X1 U1902 ( .A(n2022), .B(n225), .Y(n2023) );
  MXI2X1 U1903 ( .A(n2020), .B(n226), .S0(n432), .Y(\U3/U15/Z_4 ) );
  XNOR2X1 U1904 ( .A(n2024), .B(n2025), .Y(n2020) );
  XNOR2X1 U1905 ( .A(n2022), .B(n2019), .Y(n2025) );
  OAI21XL U1906 ( .A0(n2026), .A1(img_counter[5]), .B0(n2027), .Y(n2022) );
  OAI2BB1X1 U1907 ( .A0N(img_counter[5]), .A1N(n2026), .B0(n430), .Y(n2027) );
  XOR2X1 U1908 ( .A(n429), .B(img_counter[6]), .Y(n2024) );
  MXI2X1 U1909 ( .A(n2019), .B(n227), .S0(n432), .Y(\U3/U15/Z_3 ) );
  XNOR2X1 U1910 ( .A(n2028), .B(n2026), .Y(n2019) );
  NOR2X1 U1911 ( .A(n227), .B(n431), .Y(n2026) );
  XOR2X1 U1912 ( .A(n430), .B(img_counter[5]), .Y(n2028) );
  CLKINVX1 U1913 ( .A(n2305), .Y(\U3/U13/Z_3 ) );
  NAND2X1 U1914 ( .A(n432), .B(img_counter[3]), .Y(n2305) );
  CLKINVX1 U1915 ( .A(n2306), .Y(\U3/U13/Z_2 ) );
  NAND2X1 U1916 ( .A(n432), .B(img_counter[2]), .Y(n2306) );
  AND2X1 U1917 ( .A(N966), .B(n432), .Y(\U3/U12/Z_6 ) );
  NAND2X1 U1918 ( .A(n228), .B(n1290), .Y(\U3/U11/Z_3 ) );
  NAND2X1 U1919 ( .A(n229), .B(n1290), .Y(\U3/U11/Z_2 ) );
  NOR2X1 U1920 ( .A(n432), .B(n230), .Y(\U3/U11/Z_1 ) );
  NAND2X1 U1921 ( .A(n231), .B(n1290), .Y(\U3/U11/Z_0 ) );
  MXI2X1 U1922 ( .A(n424), .B(n230), .S0(n432), .Y(\U3/U10/Z_3 ) );
  OAI21XL U1923 ( .A0(n432), .A1(n425), .B0(n2307), .Y(\U3/U10/Z_2 ) );
  NAND2X1 U1924 ( .A(n432), .B(img_counter[0]), .Y(n2307) );
  NOR2X1 U1925 ( .A(n432), .B(n426), .Y(\U3/U10/Z_1 ) );
  NOR2X1 U1926 ( .A(n432), .B(n2029), .Y(N999) );
  XOR2X1 U1927 ( .A(n431), .B(img_counter[4]), .Y(n2029) );
endmodule

