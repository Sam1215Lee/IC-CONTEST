
module S2 ( clk, rst, S2_done, RB2_RW, RB2_A, RB2_D, RB2_Q, sen, sd );
  output [2:0] RB2_A;
  output [17:0] RB2_D;
  input [17:0] RB2_Q;
  input clk, rst, sen, sd;
  output S2_done, RB2_RW;
  wire   n168, N51, N53, N84, N85, N86, N87, N88, n6, n7, n9, n10, n11, n12,
         n13, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n151, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167;
  wire   [4:0] cnt;

  DFFSX1 \cnt_reg[2]  ( .D(n130), .CK(clk), .SN(n167), .Q(cnt[2]), .QN(n165)
         );
  DFFRX1 \cnt_reg[1]  ( .D(n114), .CK(clk), .RN(n167), .Q(cnt[1]), .QN(n6) );
  DFFRX1 \cnt_reg[0]  ( .D(n112), .CK(clk), .RN(n167), .Q(cnt[0]), .QN(n7) );
  DFFSX1 RB2_RW_reg ( .D(n107), .CK(clk), .SN(n167), .Q(n168) );
  DFFRXL \RB2_D_reg[0]  ( .D(n100), .CK(clk), .RN(n167), .QN(n95) );
  DFFRXL \RB2_D_reg[16]  ( .D(n118), .CK(clk), .RN(n167), .QN(n94) );
  DFFRXL \RB2_D_reg[12]  ( .D(n122), .CK(clk), .RN(n167), .QN(n93) );
  DFFRXL \RB2_D_reg[8]  ( .D(n111), .CK(clk), .RN(n167), .QN(n92) );
  DFFRXL \RB2_D_reg[4]  ( .D(n99), .CK(clk), .RN(n167), .QN(n91) );
  DFFRXL \RB2_D_reg[14]  ( .D(n120), .CK(clk), .RN(n167), .QN(n90) );
  DFFRXL \RB2_D_reg[10]  ( .D(n97), .CK(clk), .RN(n167), .QN(n89) );
  DFFRXL \RB2_D_reg[6]  ( .D(n98), .CK(clk), .RN(n167), .QN(n88) );
  DFFRXL \RB2_D_reg[2]  ( .D(n105), .CK(clk), .RN(n167), .QN(n87) );
  DFFRXL \RB2_D_reg[15]  ( .D(n119), .CK(clk), .RN(n167), .QN(n86) );
  DFFRXL \RB2_D_reg[11]  ( .D(n125), .CK(clk), .RN(n167), .QN(n85) );
  DFFRXL \RB2_D_reg[7]  ( .D(n109), .CK(clk), .RN(n167), .QN(n84) );
  DFFRXL \RB2_D_reg[3]  ( .D(n106), .CK(clk), .RN(n167), .QN(n83) );
  DFFRXL \RB2_D_reg[17]  ( .D(n117), .CK(clk), .RN(n167), .QN(n82) );
  DFFRXL \RB2_D_reg[13]  ( .D(n121), .CK(clk), .RN(n167), .QN(n81) );
  DFFRXL \RB2_D_reg[9]  ( .D(n110), .CK(clk), .RN(n167), .QN(n80) );
  DFFRXL \RB2_D_reg[5]  ( .D(n102), .CK(clk), .RN(n167), .QN(n79) );
  DFFRXL \RB2_D_reg[1]  ( .D(n103), .CK(clk), .RN(n167), .QN(n78) );
  DFFRXL S2_done_reg ( .D(n116), .CK(clk), .RN(n167), .QN(n77) );
  DFFRXL \RB2_A_reg[1]  ( .D(n104), .CK(clk), .RN(n167), .QN(n76) );
  DFFRXL \RB2_A_reg[2]  ( .D(n108), .CK(clk), .RN(n167), .QN(n75) );
  DFFRXL \RB2_A_reg[0]  ( .D(n101), .CK(clk), .RN(n167), .QN(n73) );
  DFFRX1 \cnt_reg[3]  ( .D(n129), .CK(clk), .RN(n167), .Q(cnt[3]) );
  DFFSX1 \cnt_reg[4]  ( .D(n127), .CK(clk), .SN(n167), .Q(cnt[4]) );
  DLY4X4 U77 ( .A(cnt[4]), .Y(n126) );
  XOR2XL U78 ( .A(n126), .B(n164), .Y(N53) );
  DLY4X4 U79 ( .A(N88), .Y(n127) );
  DLY4X1 U80 ( .A(N87), .Y(n129) );
  NOR2X6 U81 ( .A(n156), .B(n49), .Y(N87) );
  NAND2XL U82 ( .A(n162), .B(n165), .Y(n163) );
  CLKBUFX3 U83 ( .A(n6), .Y(n124) );
  OAI2BB2XL U84 ( .B0(n10), .B1(n161), .A0N(n10), .A1N(RB2_A[2]), .Y(n70) );
  OAI2BB1X1 U85 ( .A0N(RB2_RW), .A1N(n9), .B0(n10), .Y(n50) );
  NOR2X1 U86 ( .A(n113), .B(n49), .Y(N85) );
  AOI21X1 U87 ( .A0(n115), .A1(cnt[1]), .B0(n162), .Y(n157) );
  OR2X1 U88 ( .A(N51), .B(n49), .Y(N86) );
  AND2X2 U89 ( .A(sd), .B(n158), .Y(n74) );
  AO22X1 U90 ( .A0(n126), .A1(n128), .B0(n166), .B1(n126), .Y(n96) );
  DLY4X1 U91 ( .A(n59), .Y(n97) );
  DLY4X1 U92 ( .A(n63), .Y(n98) );
  DLY4X1 U93 ( .A(n65), .Y(n99) );
  DLY4X1 U94 ( .A(n69), .Y(n100) );
  DLY4X1 U95 ( .A(n72), .Y(n101) );
  NAND4BXL U96 ( .AN(n128), .B(cnt[1]), .C(n126), .D(n165), .Y(n47) );
  DLY4X1 U97 ( .A(n64), .Y(n102) );
  DLY4X1 U98 ( .A(n68), .Y(n103) );
  DLY4X1 U99 ( .A(n71), .Y(n104) );
  DLY4X1 U100 ( .A(n67), .Y(n105) );
  DLY4X1 U101 ( .A(n66), .Y(n106) );
  NAND2XL U102 ( .A(n19), .B(n39), .Y(n41) );
  DLY4X1 U103 ( .A(n50), .Y(n107) );
  DLY4X1 U104 ( .A(n70), .Y(n108) );
  NOR4BXL U105 ( .AN(n126), .B(n165), .C(n18), .D(n128), .Y(n45) );
  DLY4X1 U106 ( .A(n62), .Y(n109) );
  DLY4X1 U107 ( .A(n60), .Y(n110) );
  DLY4X1 U108 ( .A(n61), .Y(n111) );
  DLY4X1 U109 ( .A(N84), .Y(n112) );
  NOR2XL U110 ( .A(n115), .B(n49), .Y(N84) );
  DLY4X1 U111 ( .A(n157), .Y(n113) );
  DLY4X1 U112 ( .A(N85), .Y(n114) );
  DLY4X1 U113 ( .A(cnt[0]), .Y(n115) );
  DLY4X1 U114 ( .A(n51), .Y(n116) );
  DLY4X1 U115 ( .A(n52), .Y(n117) );
  DLY4X1 U116 ( .A(n53), .Y(n118) );
  NAND3BXL U117 ( .AN(n128), .B(n126), .C(n19), .Y(n15) );
  DLY4X1 U118 ( .A(n54), .Y(n119) );
  DLY4X1 U119 ( .A(n55), .Y(n120) );
  DLY4X1 U120 ( .A(n56), .Y(n121) );
  DLY4X1 U121 ( .A(n57), .Y(n122) );
  DLY4X1 U122 ( .A(n7), .Y(n123) );
  DLY4X1 U123 ( .A(n58), .Y(n125) );
  OR2XL U124 ( .A(N53), .B(n49), .Y(N88) );
  DLY4X4 U125 ( .A(cnt[3]), .Y(n128) );
  XOR2XL U126 ( .A(n128), .B(n163), .Y(n156) );
  DLY4X1 U127 ( .A(n131), .Y(n130) );
  DLY2X1 U128 ( .A(N86), .Y(n131) );
  INVX12 U129 ( .A(n77), .Y(S2_done) );
  INVX12 U130 ( .A(n82), .Y(RB2_D[17]) );
  INVX12 U131 ( .A(n94), .Y(RB2_D[16]) );
  INVX12 U132 ( .A(n86), .Y(RB2_D[15]) );
  INVX12 U133 ( .A(n90), .Y(RB2_D[14]) );
  INVX12 U134 ( .A(n81), .Y(RB2_D[13]) );
  INVX12 U135 ( .A(n93), .Y(RB2_D[12]) );
  INVX12 U136 ( .A(n85), .Y(RB2_D[11]) );
  INVX12 U137 ( .A(n89), .Y(RB2_D[10]) );
  INVX12 U138 ( .A(n80), .Y(RB2_D[9]) );
  INVX12 U139 ( .A(n92), .Y(RB2_D[8]) );
  INVX12 U140 ( .A(n84), .Y(RB2_D[7]) );
  INVX12 U141 ( .A(n88), .Y(RB2_D[6]) );
  INVX12 U142 ( .A(n79), .Y(RB2_D[5]) );
  INVX12 U143 ( .A(n91), .Y(RB2_D[4]) );
  INVX12 U144 ( .A(n83), .Y(RB2_D[3]) );
  INVX12 U145 ( .A(n87), .Y(RB2_D[2]) );
  INVX12 U146 ( .A(n78), .Y(RB2_D[1]) );
  INVX12 U147 ( .A(n95), .Y(RB2_D[0]) );
  INVXL U148 ( .A(n168), .Y(n151) );
  INVX12 U149 ( .A(n151), .Y(RB2_RW) );
  INVX12 U150 ( .A(n75), .Y(RB2_A[2]) );
  INVX12 U151 ( .A(n76), .Y(RB2_A[1]) );
  INVX12 U152 ( .A(n73), .Y(RB2_A[0]) );
  INVX6 U153 ( .A(rst), .Y(n167) );
  CLKINVX1 U154 ( .A(sen), .Y(n158) );
  NAND2X1 U155 ( .A(n123), .B(n124), .Y(n18) );
  NAND2X1 U156 ( .A(n44), .B(n158), .Y(n49) );
  AOI2BB1X1 U157 ( .A0N(n96), .A1N(n44), .B0(sen), .Y(n9) );
  CLKINVX1 U158 ( .A(n74), .Y(n161) );
  CLKINVX1 U159 ( .A(n74), .Y(n160) );
  CLKINVX1 U160 ( .A(n74), .Y(n159) );
  NAND2X1 U161 ( .A(n28), .B(n39), .Y(n35) );
  NAND2X1 U162 ( .A(n27), .B(n19), .Y(n30) );
  NAND2X1 U163 ( .A(n27), .B(n28), .Y(n21) );
  NOR2X1 U164 ( .A(sen), .B(n45), .Y(n10) );
  OAI2BB2XL U165 ( .B0(sen), .B1(n11), .A0N(S2_done), .A1N(n11), .Y(n51) );
  NOR2X1 U166 ( .A(n12), .B(sen), .Y(n11) );
  OAI2BB2XL U167 ( .B0(n43), .B1(n160), .A0N(RB2_D[1]), .A1N(n43), .Y(n68) );
  AOI2BB1X1 U168 ( .A0N(n16), .A1N(n41), .B0(sen), .Y(n43) );
  OAI2BB2XL U169 ( .B0(n37), .B1(n161), .A0N(RB2_D[5]), .A1N(n37), .Y(n64) );
  AOI2BB1X1 U170 ( .A0N(n16), .A1N(n35), .B0(sen), .Y(n37) );
  OAI2BB2XL U171 ( .B0(n32), .B1(n159), .A0N(RB2_D[9]), .A1N(n32), .Y(n60) );
  AOI2BB1X1 U172 ( .A0N(n16), .A1N(n30), .B0(sen), .Y(n32) );
  OAI2BB2XL U173 ( .B0(n25), .B1(n160), .A0N(RB2_D[13]), .A1N(n25), .Y(n56) );
  AOI2BB1X1 U174 ( .A0N(n16), .A1N(n21), .B0(sen), .Y(n25) );
  OAI2BB2XL U175 ( .B0(n13), .B1(n161), .A0N(RB2_D[17]), .A1N(n13), .Y(n52) );
  AOI2BB1X1 U176 ( .A0N(n15), .A1N(n16), .B0(sen), .Y(n13) );
  OAI2BB2XL U177 ( .B0(n40), .B1(n159), .A0N(RB2_D[3]), .A1N(n40), .Y(n66) );
  AOI2BB1X1 U178 ( .A0N(n22), .A1N(n41), .B0(sen), .Y(n40) );
  OAI2BB2XL U179 ( .B0(n34), .B1(n160), .A0N(RB2_D[7]), .A1N(n34), .Y(n62) );
  AOI2BB1X1 U180 ( .A0N(n22), .A1N(n35), .B0(sen), .Y(n34) );
  OAI2BB2XL U181 ( .B0(n29), .B1(n161), .A0N(RB2_D[11]), .A1N(n29), .Y(n58) );
  AOI2BB1X1 U182 ( .A0N(n22), .A1N(n30), .B0(sen), .Y(n29) );
  OAI2BB2XL U183 ( .B0(n20), .B1(n159), .A0N(RB2_D[15]), .A1N(n20), .Y(n54) );
  AOI2BB1X1 U184 ( .A0N(n21), .A1N(n22), .B0(sen), .Y(n20) );
  OAI2BB2XL U185 ( .B0(n42), .B1(n161), .A0N(RB2_D[2]), .A1N(n42), .Y(n67) );
  AOI2BB1X1 U186 ( .A0N(n24), .A1N(n41), .B0(sen), .Y(n42) );
  OAI2BB2XL U187 ( .B0(n36), .B1(n159), .A0N(RB2_D[6]), .A1N(n36), .Y(n63) );
  AOI2BB1X1 U188 ( .A0N(n24), .A1N(n35), .B0(sen), .Y(n36) );
  OAI2BB2XL U189 ( .B0(n31), .B1(n160), .A0N(RB2_D[10]), .A1N(n31), .Y(n59) );
  AOI2BB1X1 U190 ( .A0N(n24), .A1N(n30), .B0(sen), .Y(n31) );
  OAI2BB2XL U191 ( .B0(n23), .B1(n161), .A0N(RB2_D[14]), .A1N(n23), .Y(n55) );
  AOI2BB1X1 U192 ( .A0N(n21), .A1N(n24), .B0(sen), .Y(n23) );
  OAI2BB2XL U193 ( .B0(n38), .B1(n160), .A0N(RB2_D[4]), .A1N(n38), .Y(n65) );
  AOI2BB1X1 U194 ( .A0N(n18), .A1N(n35), .B0(sen), .Y(n38) );
  OAI2BB2XL U195 ( .B0(n33), .B1(n161), .A0N(RB2_D[8]), .A1N(n33), .Y(n61) );
  AOI2BB1X1 U196 ( .A0N(n18), .A1N(n30), .B0(sen), .Y(n33) );
  OAI2BB2XL U197 ( .B0(n26), .B1(n159), .A0N(RB2_D[12]), .A1N(n26), .Y(n57) );
  AOI2BB1X1 U198 ( .A0N(n18), .A1N(n21), .B0(sen), .Y(n26) );
  OAI2BB2XL U199 ( .B0(n17), .B1(n160), .A0N(RB2_D[16]), .A1N(n17), .Y(n53) );
  AOI2BB1X1 U200 ( .A0N(n18), .A1N(n15), .B0(sen), .Y(n17) );
  OAI2BB2XL U201 ( .B0(n9), .B1(n159), .A0N(RB2_D[0]), .A1N(n9), .Y(n69) );
  OAI2BB2XL U202 ( .B0(n48), .B1(n159), .A0N(n48), .A1N(RB2_A[0]), .Y(n72) );
  OA21XL U203 ( .A0(n115), .A1(n47), .B0(n158), .Y(n48) );
  OAI2BB2XL U204 ( .B0(n46), .B1(n160), .A0N(n46), .A1N(RB2_A[1]), .Y(n71) );
  NOR2X1 U205 ( .A(sen), .B(n12), .Y(n46) );
  NOR2X1 U206 ( .A(n96), .B(cnt[2]), .Y(n19) );
  NOR2X1 U207 ( .A(n96), .B(n165), .Y(n28) );
  NAND2X1 U208 ( .A(n115), .B(n124), .Y(n16) );
  NOR2X1 U209 ( .A(n128), .B(n126), .Y(n39) );
  NOR2BX1 U210 ( .AN(n128), .B(n126), .Y(n27) );
  NAND2X1 U211 ( .A(n115), .B(cnt[1]), .Y(n22) );
  NAND2X1 U212 ( .A(cnt[1]), .B(n123), .Y(n24) );
  NOR2X1 U213 ( .A(n123), .B(n47), .Y(n12) );
  NAND3BX1 U214 ( .AN(n18), .B(n165), .C(n39), .Y(n44) );
  NOR2X1 U215 ( .A(cnt[1]), .B(n115), .Y(n162) );
  OAI21XL U216 ( .A0(n162), .A1(n165), .B0(n163), .Y(N51) );
  NOR2X1 U217 ( .A(n128), .B(n163), .Y(n164) );
  OR2X1 U218 ( .A(cnt[1]), .B(cnt[2]), .Y(n166) );
endmodule

