
module LCD_CTRL_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2XL U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LCD_CTRL_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LCD_CTRL_DW01_add_1 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5;
  wire   [9:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(SUM[9]), .S(SUM[8]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  OAI21XL U1 ( .A0(A[2]), .A1(n3), .B0(B[2]), .Y(n4) );
  OAI2BB1X1 U2 ( .A0N(n1), .A1N(A[3]), .B0(n2), .Y(carry[4]) );
  OAI21XL U3 ( .A0(A[3]), .A1(n1), .B0(B[3]), .Y(n2) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(A[2]), .B0(n4), .Y(n1) );
  OAI2BB1X1 U5 ( .A0N(A[1]), .A1N(B[1]), .B0(n5), .Y(n3) );
  OAI211X1 U6 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n5) );
endmodule


module LCD_CTRL ( clk, reset, cmd, cmd_valid, IROM_Q, IROM_rd, IROM_A, 
        IRAM_valid, IRAM_D, IRAM_A, busy, done );
  input [3:0] cmd;
  input [7:0] IROM_Q;
  output [5:0] IROM_A;
  output [7:0] IRAM_D;
  output [5:0] IRAM_A;
  input clk, reset, cmd_valid;
  output IROM_rd, IRAM_valid, busy, done;
  wire   N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3327, N3330, N3331,
         N3333, N3334, N3338, N3339, N3340, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, cur_state,
         next_state, \img_buff[0][7] , \img_buff[0][6] , \img_buff[0][5] ,
         \img_buff[0][4] , \img_buff[0][3] , \img_buff[0][2] ,
         \img_buff[0][1] , \img_buff[0][0] , \img_buff[1][7] ,
         \img_buff[1][6] , \img_buff[1][5] , \img_buff[1][4] ,
         \img_buff[1][3] , \img_buff[1][2] , \img_buff[1][1] ,
         \img_buff[1][0] , \img_buff[2][7] , \img_buff[2][6] ,
         \img_buff[2][5] , \img_buff[2][4] , \img_buff[2][3] ,
         \img_buff[2][2] , \img_buff[2][1] , \img_buff[2][0] ,
         \img_buff[3][7] , \img_buff[3][6] , \img_buff[3][5] ,
         \img_buff[3][4] , \img_buff[3][3] , \img_buff[3][2] ,
         \img_buff[3][1] , \img_buff[3][0] , \img_buff[4][7] ,
         \img_buff[4][6] , \img_buff[4][5] , \img_buff[4][4] ,
         \img_buff[4][3] , \img_buff[4][2] , \img_buff[4][1] ,
         \img_buff[4][0] , \img_buff[5][7] , \img_buff[5][6] ,
         \img_buff[5][5] , \img_buff[5][4] , \img_buff[5][3] ,
         \img_buff[5][2] , \img_buff[5][1] , \img_buff[5][0] ,
         \img_buff[6][7] , \img_buff[6][6] , \img_buff[6][5] ,
         \img_buff[6][4] , \img_buff[6][3] , \img_buff[6][2] ,
         \img_buff[6][1] , \img_buff[6][0] , \img_buff[7][7] ,
         \img_buff[7][6] , \img_buff[7][5] , \img_buff[7][4] ,
         \img_buff[7][3] , \img_buff[7][2] , \img_buff[7][1] ,
         \img_buff[7][0] , \img_buff[8][7] , \img_buff[8][6] ,
         \img_buff[8][5] , \img_buff[8][4] , \img_buff[8][3] ,
         \img_buff[8][2] , \img_buff[8][1] , \img_buff[8][0] ,
         \img_buff[9][7] , \img_buff[9][6] , \img_buff[9][5] ,
         \img_buff[9][4] , \img_buff[9][3] , \img_buff[9][2] ,
         \img_buff[9][1] , \img_buff[9][0] , \img_buff[10][7] ,
         \img_buff[10][6] , \img_buff[10][5] , \img_buff[10][4] ,
         \img_buff[10][3] , \img_buff[10][2] , \img_buff[10][1] ,
         \img_buff[10][0] , \img_buff[11][7] , \img_buff[11][6] ,
         \img_buff[11][5] , \img_buff[11][4] , \img_buff[11][3] ,
         \img_buff[11][2] , \img_buff[11][1] , \img_buff[11][0] ,
         \img_buff[12][7] , \img_buff[12][6] , \img_buff[12][5] ,
         \img_buff[12][4] , \img_buff[12][3] , \img_buff[12][2] ,
         \img_buff[12][1] , \img_buff[12][0] , \img_buff[13][7] ,
         \img_buff[13][6] , \img_buff[13][5] , \img_buff[13][4] ,
         \img_buff[13][3] , \img_buff[13][2] , \img_buff[13][1] ,
         \img_buff[13][0] , \img_buff[14][7] , \img_buff[14][6] ,
         \img_buff[14][5] , \img_buff[14][4] , \img_buff[14][3] ,
         \img_buff[14][2] , \img_buff[14][1] , \img_buff[14][0] ,
         \img_buff[15][7] , \img_buff[15][6] , \img_buff[15][5] ,
         \img_buff[15][4] , \img_buff[15][3] , \img_buff[15][2] ,
         \img_buff[15][1] , \img_buff[15][0] , \img_buff[16][7] ,
         \img_buff[16][6] , \img_buff[16][5] , \img_buff[16][4] ,
         \img_buff[16][3] , \img_buff[16][2] , \img_buff[16][1] ,
         \img_buff[16][0] , \img_buff[17][7] , \img_buff[17][6] ,
         \img_buff[17][5] , \img_buff[17][4] , \img_buff[17][3] ,
         \img_buff[17][2] , \img_buff[17][1] , \img_buff[17][0] ,
         \img_buff[18][7] , \img_buff[18][6] , \img_buff[18][5] ,
         \img_buff[18][4] , \img_buff[18][3] , \img_buff[18][2] ,
         \img_buff[18][1] , \img_buff[18][0] , \img_buff[19][7] ,
         \img_buff[19][6] , \img_buff[19][5] , \img_buff[19][4] ,
         \img_buff[19][3] , \img_buff[19][2] , \img_buff[19][1] ,
         \img_buff[19][0] , \img_buff[20][7] , \img_buff[20][6] ,
         \img_buff[20][5] , \img_buff[20][4] , \img_buff[20][3] ,
         \img_buff[20][2] , \img_buff[20][1] , \img_buff[20][0] ,
         \img_buff[21][7] , \img_buff[21][6] , \img_buff[21][5] ,
         \img_buff[21][4] , \img_buff[21][3] , \img_buff[21][2] ,
         \img_buff[21][1] , \img_buff[21][0] , \img_buff[22][7] ,
         \img_buff[22][6] , \img_buff[22][5] , \img_buff[22][4] ,
         \img_buff[22][3] , \img_buff[22][2] , \img_buff[22][1] ,
         \img_buff[22][0] , \img_buff[23][7] , \img_buff[23][6] ,
         \img_buff[23][5] , \img_buff[23][4] , \img_buff[23][3] ,
         \img_buff[23][2] , \img_buff[23][1] , \img_buff[23][0] ,
         \img_buff[24][7] , \img_buff[24][6] , \img_buff[24][5] ,
         \img_buff[24][4] , \img_buff[24][3] , \img_buff[24][2] ,
         \img_buff[24][1] , \img_buff[24][0] , \img_buff[25][7] ,
         \img_buff[25][6] , \img_buff[25][5] , \img_buff[25][4] ,
         \img_buff[25][3] , \img_buff[25][2] , \img_buff[25][1] ,
         \img_buff[25][0] , \img_buff[26][7] , \img_buff[26][6] ,
         \img_buff[26][5] , \img_buff[26][4] , \img_buff[26][3] ,
         \img_buff[26][2] , \img_buff[26][1] , \img_buff[26][0] ,
         \img_buff[27][7] , \img_buff[27][6] , \img_buff[27][5] ,
         \img_buff[27][4] , \img_buff[27][3] , \img_buff[27][2] ,
         \img_buff[27][1] , \img_buff[27][0] , \img_buff[28][7] ,
         \img_buff[28][6] , \img_buff[28][5] , \img_buff[28][4] ,
         \img_buff[28][3] , \img_buff[28][2] , \img_buff[28][1] ,
         \img_buff[28][0] , \img_buff[29][7] , \img_buff[29][6] ,
         \img_buff[29][5] , \img_buff[29][4] , \img_buff[29][3] ,
         \img_buff[29][2] , \img_buff[29][1] , \img_buff[29][0] ,
         \img_buff[30][7] , \img_buff[30][6] , \img_buff[30][5] ,
         \img_buff[30][4] , \img_buff[30][3] , \img_buff[30][2] ,
         \img_buff[30][1] , \img_buff[30][0] , \img_buff[31][7] ,
         \img_buff[31][6] , \img_buff[31][5] , \img_buff[31][4] ,
         \img_buff[31][3] , \img_buff[31][2] , \img_buff[31][1] ,
         \img_buff[31][0] , \img_buff[32][7] , \img_buff[32][6] ,
         \img_buff[32][5] , \img_buff[32][4] , \img_buff[32][3] ,
         \img_buff[32][2] , \img_buff[32][1] , \img_buff[32][0] ,
         \img_buff[33][7] , \img_buff[33][6] , \img_buff[33][5] ,
         \img_buff[33][4] , \img_buff[33][3] , \img_buff[33][2] ,
         \img_buff[33][1] , \img_buff[33][0] , \img_buff[34][7] ,
         \img_buff[34][6] , \img_buff[34][5] , \img_buff[34][4] ,
         \img_buff[34][3] , \img_buff[34][2] , \img_buff[34][1] ,
         \img_buff[34][0] , \img_buff[35][7] , \img_buff[35][6] ,
         \img_buff[35][5] , \img_buff[35][4] , \img_buff[35][3] ,
         \img_buff[35][2] , \img_buff[35][1] , \img_buff[35][0] ,
         \img_buff[36][7] , \img_buff[36][6] , \img_buff[36][5] ,
         \img_buff[36][4] , \img_buff[36][3] , \img_buff[36][2] ,
         \img_buff[36][1] , \img_buff[36][0] , \img_buff[37][7] ,
         \img_buff[37][6] , \img_buff[37][5] , \img_buff[37][4] ,
         \img_buff[37][3] , \img_buff[37][2] , \img_buff[37][1] ,
         \img_buff[37][0] , \img_buff[38][7] , \img_buff[38][6] ,
         \img_buff[38][5] , \img_buff[38][4] , \img_buff[38][3] ,
         \img_buff[38][2] , \img_buff[38][1] , \img_buff[38][0] ,
         \img_buff[39][7] , \img_buff[39][6] , \img_buff[39][5] ,
         \img_buff[39][4] , \img_buff[39][3] , \img_buff[39][2] ,
         \img_buff[39][1] , \img_buff[39][0] , \img_buff[40][7] ,
         \img_buff[40][6] , \img_buff[40][5] , \img_buff[40][4] ,
         \img_buff[40][3] , \img_buff[40][2] , \img_buff[40][1] ,
         \img_buff[40][0] , \img_buff[41][7] , \img_buff[41][6] ,
         \img_buff[41][5] , \img_buff[41][4] , \img_buff[41][3] ,
         \img_buff[41][2] , \img_buff[41][1] , \img_buff[41][0] ,
         \img_buff[42][7] , \img_buff[42][6] , \img_buff[42][5] ,
         \img_buff[42][4] , \img_buff[42][3] , \img_buff[42][2] ,
         \img_buff[42][1] , \img_buff[42][0] , \img_buff[43][7] ,
         \img_buff[43][6] , \img_buff[43][5] , \img_buff[43][4] ,
         \img_buff[43][3] , \img_buff[43][2] , \img_buff[43][1] ,
         \img_buff[43][0] , \img_buff[44][7] , \img_buff[44][6] ,
         \img_buff[44][5] , \img_buff[44][4] , \img_buff[44][3] ,
         \img_buff[44][2] , \img_buff[44][1] , \img_buff[44][0] ,
         \img_buff[45][7] , \img_buff[45][6] , \img_buff[45][5] ,
         \img_buff[45][4] , \img_buff[45][3] , \img_buff[45][2] ,
         \img_buff[45][1] , \img_buff[45][0] , \img_buff[46][7] ,
         \img_buff[46][6] , \img_buff[46][5] , \img_buff[46][4] ,
         \img_buff[46][3] , \img_buff[46][2] , \img_buff[46][1] ,
         \img_buff[46][0] , \img_buff[47][7] , \img_buff[47][6] ,
         \img_buff[47][5] , \img_buff[47][4] , \img_buff[47][3] ,
         \img_buff[47][2] , \img_buff[47][1] , \img_buff[47][0] ,
         \img_buff[48][7] , \img_buff[48][6] , \img_buff[48][5] ,
         \img_buff[48][4] , \img_buff[48][3] , \img_buff[48][2] ,
         \img_buff[48][1] , \img_buff[48][0] , \img_buff[49][7] ,
         \img_buff[49][6] , \img_buff[49][5] , \img_buff[49][4] ,
         \img_buff[49][3] , \img_buff[49][2] , \img_buff[49][1] ,
         \img_buff[49][0] , \img_buff[50][7] , \img_buff[50][6] ,
         \img_buff[50][5] , \img_buff[50][4] , \img_buff[50][3] ,
         \img_buff[50][2] , \img_buff[50][1] , \img_buff[50][0] ,
         \img_buff[51][7] , \img_buff[51][6] , \img_buff[51][5] ,
         \img_buff[51][4] , \img_buff[51][3] , \img_buff[51][2] ,
         \img_buff[51][1] , \img_buff[51][0] , \img_buff[52][7] ,
         \img_buff[52][6] , \img_buff[52][5] , \img_buff[52][4] ,
         \img_buff[52][3] , \img_buff[52][2] , \img_buff[52][1] ,
         \img_buff[52][0] , \img_buff[53][7] , \img_buff[53][6] ,
         \img_buff[53][5] , \img_buff[53][4] , \img_buff[53][3] ,
         \img_buff[53][2] , \img_buff[53][1] , \img_buff[53][0] ,
         \img_buff[54][7] , \img_buff[54][6] , \img_buff[54][5] ,
         \img_buff[54][4] , \img_buff[54][3] , \img_buff[54][2] ,
         \img_buff[54][1] , \img_buff[54][0] , \img_buff[55][7] ,
         \img_buff[55][6] , \img_buff[55][5] , \img_buff[55][4] ,
         \img_buff[55][3] , \img_buff[55][2] , \img_buff[55][1] ,
         \img_buff[55][0] , \img_buff[56][7] , \img_buff[56][6] ,
         \img_buff[56][5] , \img_buff[56][4] , \img_buff[56][3] ,
         \img_buff[56][2] , \img_buff[56][1] , \img_buff[56][0] ,
         \img_buff[57][7] , \img_buff[57][6] , \img_buff[57][5] ,
         \img_buff[57][4] , \img_buff[57][3] , \img_buff[57][2] ,
         \img_buff[57][1] , \img_buff[57][0] , \img_buff[58][7] ,
         \img_buff[58][6] , \img_buff[58][5] , \img_buff[58][4] ,
         \img_buff[58][3] , \img_buff[58][2] , \img_buff[58][1] ,
         \img_buff[58][0] , \img_buff[59][7] , \img_buff[59][6] ,
         \img_buff[59][5] , \img_buff[59][4] , \img_buff[59][3] ,
         \img_buff[59][2] , \img_buff[59][1] , \img_buff[59][0] ,
         \img_buff[60][7] , \img_buff[60][6] , \img_buff[60][5] ,
         \img_buff[60][4] , \img_buff[60][3] , \img_buff[60][2] ,
         \img_buff[60][1] , \img_buff[60][0] , \img_buff[61][7] ,
         \img_buff[61][6] , \img_buff[61][5] , \img_buff[61][4] ,
         \img_buff[61][3] , \img_buff[61][2] , \img_buff[61][1] ,
         \img_buff[61][0] , \img_buff[62][7] , \img_buff[62][6] ,
         \img_buff[62][5] , \img_buff[62][4] , \img_buff[62][3] ,
         \img_buff[62][2] , \img_buff[62][1] , \img_buff[62][0] ,
         \img_buff[63][7] , \img_buff[63][6] , \img_buff[63][5] ,
         \img_buff[63][4] , \img_buff[63][3] , \img_buff[63][2] ,
         \img_buff[63][1] , \img_buff[63][0] , N3344, N3345, N3346, N3347,
         N3348, N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3357, N3358,
         N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3369,
         N3375, N3380, N3381, N3382, N3383, N3384, N3385, N3451, N3452, N3453,
         N3454, N3455, N3490, N3491, N3492, N4817, N4818, N4819, N5079, N5080,
         N5081, N5341, N5342, N5343, N5602, N5603, N5604, N6161, N6162, N6163,
         N6164, N6165, N6166, N16287, n93, n162, n164, n166, n168, n170, n172,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n944, n963,
         n964, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n982, n983, n984, n985, n986, n989,
         n991, n993, n994, n996, n997, n998, n999, n1001, n1002, n1003, n1004,
         n1006, n1007, n1008, n1009, n1011, n1012, n1013, n1014, n1016, n1017,
         n1018, n1019, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1096, n1097, n1098, n1099, n1100,
         n1102, n1104, n1105, n1106, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1116, n1117, n1118, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1132, n1133, n1134, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, N6160, N6159, N6158, N6157, N6156, N6155, N6154, N6153, N6152,
         N6151, N6150, N6149, N6148, N6147, N6146, N6145, N6144, N6143,
         \add_139/carry[5] , \add_139/carry[4] , \add_139/carry[3] ,
         \add_139/carry[2] , \add_118/carry[5] , \add_118/carry[4] ,
         \add_118/carry[3] , \add_118/carry[2] , \sub_80/carry[2] ,
         \sub_80/carry[3] , n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4729, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666;
  wire   [3:0] cmd_reg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign done = 1'b1;

  DFFRX4 cur_state_reg ( .D(next_state), .CK(clk), .RN(n6642), .Q(cur_state), 
        .QN(n93) );
  AOI221X2 U63 ( .A0(n4701), .A1(n1023), .B0(n4697), .B1(n1045), .C0(n1046), 
        .Y(n1039) );
  OAI221X2 U67 ( .A0(n5779), .A1(n1025), .B0(n4658), .B1(n1027), .C0(n1056), 
        .Y(n1045) );
  AOI221X2 U525 ( .A0(n1498), .A1(n4701), .B0(n4697), .B1(n1512), .C0(n1513), 
        .Y(n1510) );
  OAI221X2 U529 ( .A0(n5777), .A1(n1500), .B0(n4663), .B1(n1507), .C0(n1516), 
        .Y(n1512) );
  AOI221X2 U572 ( .A0(n1542), .A1(n4701), .B0(n4697), .B1(n1556), .C0(n1557), 
        .Y(n1554) );
  OAI221X2 U576 ( .A0(n5777), .A1(n1544), .B0(n4664), .B1(n1551), .C0(n1560), 
        .Y(n1556) );
  AOI221X2 U619 ( .A0(n1586), .A1(n4701), .B0(n4697), .B1(n1600), .C0(n1601), 
        .Y(n1598) );
  OAI22X4 U667 ( .A0(n5913), .A1(n1633), .B0(n1646), .B1(n4637), .Y(n1645) );
  OAI22X4 U714 ( .A0(n5913), .A1(n1677), .B0(n1690), .B1(n4637), .Y(n1689) );
  OAI22X4 U761 ( .A0(n5913), .A1(n1721), .B0(n1734), .B1(n4637), .Y(n1733) );
  AOI221X2 U808 ( .A0(n1762), .A1(n4701), .B0(n4697), .B1(n1777), .C0(n1778), 
        .Y(n1774) );
  AOI221X2 U859 ( .A0(n1807), .A1(n4701), .B0(n4697), .B1(n1821), .C0(n1822), 
        .Y(n1819) );
  AOI221X2 U906 ( .A0(n1851), .A1(n4701), .B0(n4697), .B1(n1864), .C0(n1865), 
        .Y(n1863) );
  AOI221X2 U953 ( .A0(n1890), .A1(n4701), .B0(n4697), .B1(n1903), .C0(n1904), 
        .Y(n1902) );
  OAI22X4 U954 ( .A0(n5913), .A1(n1893), .B0(n1905), .B1(n4637), .Y(n1904) );
  AOI221X2 U1000 ( .A0(n1929), .A1(n4701), .B0(n4697), .B1(n1942), .C0(n1943), 
        .Y(n1941) );
  AOI221X2 U1047 ( .A0(n1968), .A1(n4701), .B0(n4697), .B1(n1981), .C0(n1982), 
        .Y(n1980) );
  OAI22X4 U1048 ( .A0(n5913), .A1(n1971), .B0(n1983), .B1(n4637), .Y(n1982) );
  AOI221X2 U1094 ( .A0(n2007), .A1(n4701), .B0(n4697), .B1(n2021), .C0(n2022), 
        .Y(n2020) );
  AOI221X2 U1141 ( .A0(n2048), .A1(n4701), .B0(n4697), .B1(n2059), .C0(n2060), 
        .Y(n2058) );
  OAI22X4 U1142 ( .A0(n5914), .A1(n2051), .B0(n2061), .B1(n4637), .Y(n2060) );
  AOI221X2 U1189 ( .A0(n2087), .A1(n4701), .B0(n4697), .B1(n2098), .C0(n2099), 
        .Y(n2097) );
  OAI22X4 U1190 ( .A0(n5914), .A1(n2090), .B0(n2100), .B1(n4637), .Y(n2099) );
  AOI221X2 U1240 ( .A0(n2126), .A1(n4701), .B0(n4697), .B1(n2138), .C0(n2139), 
        .Y(n2136) );
  OAI22X4 U1241 ( .A0(n5914), .A1(n2129), .B0(n2140), .B1(n4637), .Y(n2139) );
  AOI221X2 U1287 ( .A0(n2170), .A1(n4701), .B0(n4697), .B1(n2181), .C0(n2182), 
        .Y(n2180) );
  OAI22X4 U1288 ( .A0(n5914), .A1(n2173), .B0(n2183), .B1(n4637), .Y(n2182) );
  AOI221X2 U1334 ( .A0(n2209), .A1(n4701), .B0(n4697), .B1(n2220), .C0(n2221), 
        .Y(n2219) );
  OAI22X4 U1335 ( .A0(n5914), .A1(n2212), .B0(n2222), .B1(n4637), .Y(n2221) );
  AOI221X2 U1381 ( .A0(n2248), .A1(n4701), .B0(n4697), .B1(n2259), .C0(n2260), 
        .Y(n2258) );
  OAI22X4 U1382 ( .A0(n5914), .A1(n2251), .B0(n2261), .B1(n4637), .Y(n2260) );
  AOI221X2 U1428 ( .A0(n2287), .A1(n4701), .B0(n4697), .B1(n2298), .C0(n2299), 
        .Y(n2297) );
  OAI22X4 U1429 ( .A0(n5914), .A1(n2290), .B0(n2300), .B1(n4637), .Y(n2299) );
  AOI221X2 U1475 ( .A0(n2326), .A1(n4701), .B0(n4697), .B1(n2337), .C0(n2338), 
        .Y(n2336) );
  OAI22X4 U1476 ( .A0(n5914), .A1(n2329), .B0(n2339), .B1(n4637), .Y(n2338) );
  AOI221X2 U1522 ( .A0(n2365), .A1(n4701), .B0(n4697), .B1(n2376), .C0(n2377), 
        .Y(n2375) );
  OAI22X4 U1523 ( .A0(n5914), .A1(n2368), .B0(n2378), .B1(n4637), .Y(n2377) );
  AOI221X2 U1570 ( .A0(n2404), .A1(n4701), .B0(n4697), .B1(n2415), .C0(n2416), 
        .Y(n2414) );
  OAI22X4 U1571 ( .A0(n5914), .A1(n2407), .B0(n2417), .B1(n4637), .Y(n2416) );
  AOI221X2 U1621 ( .A0(n2443), .A1(n4701), .B0(n4697), .B1(n2455), .C0(n2456), 
        .Y(n2453) );
  OAI22X4 U1622 ( .A0(n5914), .A1(n2446), .B0(n2457), .B1(n4637), .Y(n2456) );
  AOI221X2 U1668 ( .A0(n2487), .A1(n4701), .B0(n4697), .B1(n2498), .C0(n2499), 
        .Y(n2497) );
  OAI22X4 U1669 ( .A0(n5914), .A1(n2490), .B0(n2500), .B1(n4637), .Y(n2499) );
  AOI221X2 U1670 ( .A0(n6627), .A1(n4696), .B0(n6562), .B1(n4650), .C0(n2501), 
        .Y(n2500) );
  AOI221X2 U1715 ( .A0(n2526), .A1(n4701), .B0(n4697), .B1(n2537), .C0(n2538), 
        .Y(n2536) );
  OAI22X4 U1716 ( .A0(n5914), .A1(n2529), .B0(n2539), .B1(n4637), .Y(n2538) );
  AOI221X2 U1717 ( .A0(n6619), .A1(n4696), .B0(n6554), .B1(n4650), .C0(n2540), 
        .Y(n2539) );
  AOI221X2 U1762 ( .A0(n2565), .A1(n4701), .B0(n4697), .B1(n2576), .C0(n2577), 
        .Y(n2575) );
  OAI22X4 U1763 ( .A0(n5914), .A1(n2568), .B0(n2578), .B1(n4637), .Y(n2577) );
  AOI221X2 U1764 ( .A0(n6611), .A1(n4696), .B0(n6546), .B1(n4650), .C0(n2579), 
        .Y(n2578) );
  AOI221X2 U1856 ( .A0(n2643), .A1(n4701), .B0(n4697), .B1(n2654), .C0(n2655), 
        .Y(n2653) );
  OAI22X4 U1857 ( .A0(n5915), .A1(n2646), .B0(n2656), .B1(n4637), .Y(n2655) );
  AOI221X2 U1858 ( .A0(n6595), .A1(n4696), .B0(n6530), .B1(n4650), .C0(n2657), 
        .Y(n2656) );
  AOI221X2 U1951 ( .A0(n2721), .A1(n4701), .B0(n4697), .B1(n2732), .C0(n2733), 
        .Y(n2731) );
  OAI22X4 U1952 ( .A0(n5915), .A1(n2724), .B0(n2734), .B1(n4637), .Y(n2733) );
  AOI221X2 U2002 ( .A0(n2760), .A1(n4701), .B0(n4697), .B1(n2772), .C0(n2773), 
        .Y(n2770) );
  OAI22X4 U2003 ( .A0(n5915), .A1(n2763), .B0(n2774), .B1(n4637), .Y(n2773) );
  AOI221X2 U2049 ( .A0(n2804), .A1(n4701), .B0(n4697), .B1(n2815), .C0(n2816), 
        .Y(n2814) );
  OAI22X4 U2050 ( .A0(n5915), .A1(n2807), .B0(n2817), .B1(n4637), .Y(n2816) );
  AOI221X2 U2096 ( .A0(n2843), .A1(n4701), .B0(n4697), .B1(n2854), .C0(n2855), 
        .Y(n2853) );
  OAI22X4 U2097 ( .A0(n5915), .A1(n2846), .B0(n2856), .B1(n4637), .Y(n2855) );
  AOI221X2 U2143 ( .A0(n2882), .A1(n4701), .B0(n4697), .B1(n2893), .C0(n2894), 
        .Y(n2892) );
  OAI22X4 U2144 ( .A0(n5915), .A1(n2885), .B0(n2895), .B1(n4637), .Y(n2894) );
  AOI221X2 U2190 ( .A0(n2921), .A1(n4701), .B0(n4697), .B1(n2932), .C0(n2933), 
        .Y(n2931) );
  AOI221X2 U2237 ( .A0(n2960), .A1(n4701), .B0(n4697), .B1(n2971), .C0(n2972), 
        .Y(n2970) );
  OAI22X4 U2238 ( .A0(n5915), .A1(n2963), .B0(n2973), .B1(n4637), .Y(n2972) );
  AOI221X2 U2284 ( .A0(n2999), .A1(n4701), .B0(n4697), .B1(n3010), .C0(n3011), 
        .Y(n3009) );
  OAI22X4 U2285 ( .A0(n5915), .A1(n3002), .B0(n3012), .B1(n4637), .Y(n3011) );
  AOI221X2 U2332 ( .A0(n3038), .A1(n4701), .B0(n4697), .B1(n3049), .C0(n3050), 
        .Y(n3048) );
  OAI22X4 U2333 ( .A0(n5915), .A1(n3041), .B0(n3051), .B1(n4637), .Y(n3050) );
  AOI221X2 U2383 ( .A0(n3077), .A1(n4701), .B0(n4697), .B1(n3089), .C0(n3090), 
        .Y(n3087) );
  OAI22X4 U2384 ( .A0(n5915), .A1(n3080), .B0(n3091), .B1(n4637), .Y(n3090) );
  AOI221X2 U2385 ( .A0(n6633), .A1(n4696), .B0(n6568), .B1(n4650), .C0(n3092), 
        .Y(n3091) );
  AOI221X2 U2430 ( .A0(n3121), .A1(n4701), .B0(n4697), .B1(n3132), .C0(n3133), 
        .Y(n3131) );
  OAI22X4 U2431 ( .A0(n5915), .A1(n3124), .B0(n3134), .B1(n4637), .Y(n3133) );
  AOI221X2 U2432 ( .A0(n6625), .A1(n4696), .B0(n6560), .B1(n4650), .C0(n3135), 
        .Y(n3134) );
  AOI221X2 U2477 ( .A0(n3160), .A1(n4701), .B0(n4697), .B1(n3171), .C0(n3172), 
        .Y(n3170) );
  OAI22X4 U2478 ( .A0(n5915), .A1(n3163), .B0(n3173), .B1(n4637), .Y(n3172) );
  AOI221X2 U2524 ( .A0(n3199), .A1(n4701), .B0(n4697), .B1(n3210), .C0(n3211), 
        .Y(n3209) );
  AOI221X2 U2571 ( .A0(n3238), .A1(n4701), .B0(n4697), .B1(n3249), .C0(n3250), 
        .Y(n3248) );
  AOI221X2 U2618 ( .A0(n3277), .A1(n4701), .B0(n4697), .B1(n3288), .C0(n3289), 
        .Y(n3287) );
  AOI221X2 U2665 ( .A0(n3316), .A1(n4701), .B0(n4697), .B1(n3327), .C0(n3328), 
        .Y(n3326) );
  AOI221X2 U2713 ( .A0(n3355), .A1(n4701), .B0(n4697), .B1(n3366), .C0(n3367), 
        .Y(n3365) );
  AOI221X2 U2764 ( .A0(n3394), .A1(n4701), .B0(n4697), .B1(n3406), .C0(n3407), 
        .Y(n3404) );
  AOI221X2 U2811 ( .A0(n3438), .A1(n4701), .B0(n4697), .B1(n3449), .C0(n3450), 
        .Y(n3448) );
  AOI221X2 U2858 ( .A0(n3477), .A1(n4701), .B0(n4697), .B1(n3488), .C0(n3489), 
        .Y(n3487) );
  AOI221X2 U2905 ( .A0(n3516), .A1(n4701), .B0(n4697), .B1(n3527), .C0(n3528), 
        .Y(n3526) );
  OAI22X4 U2906 ( .A0(n5912), .A1(n3519), .B0(n3529), .B1(n4637), .Y(n3528) );
  AOI221X2 U3094 ( .A0(n3672), .A1(n4701), .B0(n4697), .B1(n3683), .C0(n3684), 
        .Y(n3682) );
  AOI221X2 U3250 ( .A0(n3794), .A1(n4701), .B0(n4697), .B1(n3805), .C0(n3806), 
        .Y(n3804) );
  AOI221X2 U3302 ( .A0(n3833), .A1(n4701), .B0(n4697), .B1(n3844), .C0(n3845), 
        .Y(n3843) );
  AOI221X2 U3354 ( .A0(n3872), .A1(n4701), .B0(n4697), .B1(n3883), .C0(n3884), 
        .Y(n3882) );
  AOI221X2 U3406 ( .A0(n3911), .A1(n4701), .B0(n4697), .B1(n3922), .C0(n3923), 
        .Y(n3921) );
  AOI221X2 U3459 ( .A0(n3950), .A1(n4701), .B0(n4697), .B1(n3962), .C0(n3963), 
        .Y(n3960) );
  OAI222X2 U3523 ( .A0(n4017), .A1(n3975), .B0(n4018), .B1(n5668), .C0(n4000), 
        .C1(n168), .Y(n1012) );
  AOI221X2 U3567 ( .A0(n4038), .A1(n4701), .B0(n4697), .B1(n4049), .C0(n4050), 
        .Y(n4048) );
  OAI31X2 U3671 ( .A0(n93), .A1(n4061), .A2(n1476), .B0(n6642), .Y(n4094) );
  LCD_CTRL_DW01_add_3 add_248_2 ( .A({1'b0, N3360, n5660, n5661, n5662, n5663, 
        n5664, n5665, n5666}), .B({1'b0, n5948, n5945, n5940, n5934, n5928, 
        n5925, n5920, n5918}), .CI(1'b0), .SUM({N6160, N6159, N6158, N6157, 
        N6156, N6155, N6154, N6153, N6152}) );
  LCD_CTRL_DW01_add_2 add_248 ( .A({1'b0, n5651, n5652, n5653, n5654, n5655, 
        n5656, n5657, N3351}), .B({1'b0, n5658, N3353, n5659, N3355, n4667, 
        N3357, N3358, N3359}), .CI(1'b0), .SUM({N6151, N6150, N6149, N6148, 
        N6147, N6146, N6145, N6144, N6143}) );
  LCD_CTRL_DW01_add_1 add_248_3 ( .A({1'b0, N6151, N6150, N6149, N6148, N6147, 
        N6146, N6145, N6144, N6143}), .B({1'b0, N6160, N6159, N6158, N6157, 
        N6156, N6155, N6154, N6153, N6152}), .CI(1'b0), .SUM({N6166, N6165, 
        N6164, N6163, N6162, N6161, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3}) );
  EDFFX1 \avg_reg[3]  ( .D(N6162), .E(N16287), .CK(clk), .QN(n170) );
  EDFFX1 \avg_reg[2]  ( .D(N6161), .E(N16287), .CK(clk), .QN(n172) );
  EDFFX1 \cmd_reg_reg[0]  ( .D(cmd[0]), .E(n4883), .CK(clk), .Q(cmd_reg[0]), 
        .QN(n964) );
  EDFFX1 \cmd_reg_reg[1]  ( .D(cmd[1]), .E(n4883), .CK(clk), .Q(cmd_reg[1]), 
        .QN(n963) );
  DFFX1 \img_buff_reg[1][7]  ( .D(n4104), .CK(clk), .Q(\img_buff[1][7] ), .QN(
        n206) );
  DFFX1 \img_buff_reg[5][7]  ( .D(n4136), .CK(clk), .Q(\img_buff[5][7] ), .QN(
        n238) );
  DFFX1 \img_buff_reg[9][7]  ( .D(n4168), .CK(clk), .Q(\img_buff[9][7] ), .QN(
        n270) );
  DFFX1 \img_buff_reg[13][7]  ( .D(n4200), .CK(clk), .Q(\img_buff[13][7] ), 
        .QN(n302) );
  DFFX1 \img_buff_reg[17][7]  ( .D(n4232), .CK(clk), .Q(\img_buff[17][7] ), 
        .QN(n334) );
  DFFX1 \img_buff_reg[25][7]  ( .D(n4296), .CK(clk), .Q(\img_buff[25][7] ), 
        .QN(n398) );
  DFFX1 \img_buff_reg[33][7]  ( .D(n4360), .CK(clk), .Q(\img_buff[33][7] ), 
        .QN(n462) );
  DFFX1 \img_buff_reg[37][7]  ( .D(n4392), .CK(clk), .Q(\img_buff[37][7] ), 
        .QN(n494) );
  DFFX1 \img_buff_reg[41][7]  ( .D(n4424), .CK(clk), .Q(\img_buff[41][7] ), 
        .QN(n526) );
  DFFX1 \img_buff_reg[45][7]  ( .D(n4456), .CK(clk), .Q(\img_buff[45][7] ), 
        .QN(n558) );
  DFFX1 \img_buff_reg[49][7]  ( .D(n4488), .CK(clk), .Q(\img_buff[49][7] ), 
        .QN(n590) );
  DFFX1 \img_buff_reg[57][7]  ( .D(n4552), .CK(clk), .Q(\img_buff[57][7] ), 
        .QN(n654) );
  DFFX1 \img_buff_reg[3][7]  ( .D(n4120), .CK(clk), .Q(\img_buff[3][7] ), .QN(
        n222) );
  DFFX1 \img_buff_reg[11][7]  ( .D(n4184), .CK(clk), .Q(\img_buff[11][7] ), 
        .QN(n286) );
  DFFX1 \img_buff_reg[35][7]  ( .D(n4376), .CK(clk), .Q(\img_buff[35][7] ), 
        .QN(n478) );
  DFFX1 \img_buff_reg[43][7]  ( .D(n4440), .CK(clk), .Q(\img_buff[43][7] ), 
        .QN(n542) );
  DFFX1 \img_buff_reg[4][7]  ( .D(n4128), .CK(clk), .Q(\img_buff[4][7] ), .QN(
        n230) );
  DFFX1 \img_buff_reg[8][7]  ( .D(n4160), .CK(clk), .Q(\img_buff[8][7] ), .QN(
        n262) );
  DFFX1 \img_buff_reg[12][7]  ( .D(n4192), .CK(clk), .Q(\img_buff[12][7] ), 
        .QN(n294) );
  DFFX1 \img_buff_reg[16][7]  ( .D(n4224), .CK(clk), .Q(\img_buff[16][7] ), 
        .QN(n326) );
  DFFX1 \img_buff_reg[24][7]  ( .D(n4288), .CK(clk), .Q(\img_buff[24][7] ), 
        .QN(n390) );
  DFFX1 \img_buff_reg[32][7]  ( .D(n4352), .CK(clk), .Q(\img_buff[32][7] ), 
        .QN(n454) );
  DFFX1 \img_buff_reg[36][7]  ( .D(n4384), .CK(clk), .Q(\img_buff[36][7] ), 
        .QN(n486) );
  DFFX1 \img_buff_reg[40][7]  ( .D(n4416), .CK(clk), .Q(\img_buff[40][7] ), 
        .QN(n518) );
  DFFX1 \img_buff_reg[44][7]  ( .D(n4448), .CK(clk), .Q(\img_buff[44][7] ), 
        .QN(n550) );
  DFFX1 \img_buff_reg[48][7]  ( .D(n4480), .CK(clk), .Q(\img_buff[48][7] ), 
        .QN(n582) );
  DFFX1 \img_buff_reg[56][7]  ( .D(n4544), .CK(clk), .Q(\img_buff[56][7] ), 
        .QN(n646) );
  DFFX1 \img_buff_reg[2][7]  ( .D(n4112), .CK(clk), .Q(\img_buff[2][7] ), .QN(
        n214) );
  DFFX1 \img_buff_reg[10][7]  ( .D(n4176), .CK(clk), .Q(\img_buff[10][7] ), 
        .QN(n278) );
  DFFX1 \img_buff_reg[34][7]  ( .D(n4368), .CK(clk), .Q(\img_buff[34][7] ), 
        .QN(n470) );
  DFFX1 \img_buff_reg[42][7]  ( .D(n4432), .CK(clk), .Q(\img_buff[42][7] ), 
        .QN(n534) );
  DFFX1 \img_buff_reg[1][6]  ( .D(n4105), .CK(clk), .Q(\img_buff[1][6] ), .QN(
        n207) );
  DFFX1 \img_buff_reg[5][6]  ( .D(n4137), .CK(clk), .Q(\img_buff[5][6] ), .QN(
        n239) );
  DFFX1 \img_buff_reg[9][6]  ( .D(n4169), .CK(clk), .Q(\img_buff[9][6] ), .QN(
        n271) );
  DFFX1 \img_buff_reg[13][6]  ( .D(n4201), .CK(clk), .Q(\img_buff[13][6] ), 
        .QN(n303) );
  DFFX1 \img_buff_reg[17][6]  ( .D(n4233), .CK(clk), .Q(\img_buff[17][6] ), 
        .QN(n335) );
  DFFX1 \img_buff_reg[21][6]  ( .D(n4265), .CK(clk), .Q(\img_buff[21][6] ), 
        .QN(n367) );
  DFFX1 \img_buff_reg[25][6]  ( .D(n4297), .CK(clk), .Q(\img_buff[25][6] ), 
        .QN(n399) );
  DFFX1 \img_buff_reg[29][6]  ( .D(n4329), .CK(clk), .Q(\img_buff[29][6] ), 
        .QN(n431) );
  DFFX1 \img_buff_reg[33][6]  ( .D(n4361), .CK(clk), .Q(\img_buff[33][6] ), 
        .QN(n463) );
  DFFX1 \img_buff_reg[37][6]  ( .D(n4393), .CK(clk), .Q(\img_buff[37][6] ), 
        .QN(n495) );
  DFFX1 \img_buff_reg[41][6]  ( .D(n4425), .CK(clk), .Q(\img_buff[41][6] ), 
        .QN(n527) );
  DFFX1 \img_buff_reg[45][6]  ( .D(n4457), .CK(clk), .Q(\img_buff[45][6] ), 
        .QN(n559) );
  DFFX1 \img_buff_reg[49][6]  ( .D(n4489), .CK(clk), .Q(\img_buff[49][6] ), 
        .QN(n591) );
  DFFX1 \img_buff_reg[53][6]  ( .D(n4521), .CK(clk), .Q(\img_buff[53][6] ), 
        .QN(n623) );
  DFFX1 \img_buff_reg[57][6]  ( .D(n4553), .CK(clk), .Q(\img_buff[57][6] ), 
        .QN(n655) );
  DFFX1 \img_buff_reg[61][6]  ( .D(n4585), .CK(clk), .Q(\img_buff[61][6] ), 
        .QN(n687) );
  DFFX1 \img_buff_reg[21][7]  ( .D(n4264), .CK(clk), .Q(\img_buff[21][7] ), 
        .QN(n366) );
  DFFX1 \img_buff_reg[29][7]  ( .D(n4328), .CK(clk), .Q(\img_buff[29][7] ), 
        .QN(n430) );
  DFFX1 \img_buff_reg[53][7]  ( .D(n4520), .CK(clk), .Q(\img_buff[53][7] ), 
        .QN(n622) );
  DFFX1 \img_buff_reg[61][7]  ( .D(n4584), .CK(clk), .Q(\img_buff[61][7] ), 
        .QN(n686) );
  DFFX1 \img_buff_reg[1][5]  ( .D(n4106), .CK(clk), .Q(\img_buff[1][5] ), .QN(
        n208) );
  DFFX1 \img_buff_reg[5][5]  ( .D(n4138), .CK(clk), .Q(\img_buff[5][5] ), .QN(
        n240) );
  DFFX1 \img_buff_reg[9][5]  ( .D(n4170), .CK(clk), .Q(\img_buff[9][5] ), .QN(
        n272) );
  DFFX1 \img_buff_reg[13][5]  ( .D(n4202), .CK(clk), .Q(\img_buff[13][5] ), 
        .QN(n304) );
  DFFX1 \img_buff_reg[17][5]  ( .D(n4234), .CK(clk), .Q(\img_buff[17][5] ), 
        .QN(n336) );
  DFFX1 \img_buff_reg[21][5]  ( .D(n4266), .CK(clk), .Q(\img_buff[21][5] ), 
        .QN(n368) );
  DFFX1 \img_buff_reg[25][5]  ( .D(n4298), .CK(clk), .Q(\img_buff[25][5] ), 
        .QN(n400) );
  DFFX1 \img_buff_reg[29][5]  ( .D(n4330), .CK(clk), .Q(\img_buff[29][5] ), 
        .QN(n432) );
  DFFX1 \img_buff_reg[33][5]  ( .D(n4362), .CK(clk), .Q(\img_buff[33][5] ), 
        .QN(n464) );
  DFFX1 \img_buff_reg[37][5]  ( .D(n4394), .CK(clk), .Q(\img_buff[37][5] ), 
        .QN(n496) );
  DFFX1 \img_buff_reg[41][5]  ( .D(n4426), .CK(clk), .Q(\img_buff[41][5] ), 
        .QN(n528) );
  DFFX1 \img_buff_reg[45][5]  ( .D(n4458), .CK(clk), .Q(\img_buff[45][5] ), 
        .QN(n560) );
  DFFX1 \img_buff_reg[49][5]  ( .D(n4490), .CK(clk), .Q(\img_buff[49][5] ), 
        .QN(n592) );
  DFFX1 \img_buff_reg[53][5]  ( .D(n4522), .CK(clk), .Q(\img_buff[53][5] ), 
        .QN(n624) );
  DFFX1 \img_buff_reg[57][5]  ( .D(n4554), .CK(clk), .Q(\img_buff[57][5] ), 
        .QN(n656) );
  DFFX1 \img_buff_reg[61][5]  ( .D(n4586), .CK(clk), .Q(\img_buff[61][5] ), 
        .QN(n688) );
  DFFX1 \img_buff_reg[1][3]  ( .D(n4108), .CK(clk), .Q(\img_buff[1][3] ), .QN(
        n210) );
  DFFX1 \img_buff_reg[5][3]  ( .D(n4140), .CK(clk), .Q(\img_buff[5][3] ), .QN(
        n242) );
  DFFX1 \img_buff_reg[9][3]  ( .D(n4172), .CK(clk), .Q(\img_buff[9][3] ), .QN(
        n274) );
  DFFX1 \img_buff_reg[13][3]  ( .D(n4204), .CK(clk), .Q(\img_buff[13][3] ), 
        .QN(n306) );
  DFFX1 \img_buff_reg[17][3]  ( .D(n4236), .CK(clk), .Q(\img_buff[17][3] ), 
        .QN(n338) );
  DFFX1 \img_buff_reg[21][3]  ( .D(n4268), .CK(clk), .Q(\img_buff[21][3] ), 
        .QN(n370) );
  DFFX1 \img_buff_reg[25][3]  ( .D(n4300), .CK(clk), .Q(\img_buff[25][3] ), 
        .QN(n402) );
  DFFX1 \img_buff_reg[29][3]  ( .D(n4332), .CK(clk), .Q(\img_buff[29][3] ), 
        .QN(n434) );
  DFFX1 \img_buff_reg[33][3]  ( .D(n4364), .CK(clk), .Q(\img_buff[33][3] ), 
        .QN(n466) );
  DFFX1 \img_buff_reg[37][3]  ( .D(n4396), .CK(clk), .Q(\img_buff[37][3] ), 
        .QN(n498) );
  DFFX1 \img_buff_reg[41][3]  ( .D(n4428), .CK(clk), .Q(\img_buff[41][3] ), 
        .QN(n530) );
  DFFX1 \img_buff_reg[45][3]  ( .D(n4460), .CK(clk), .Q(\img_buff[45][3] ), 
        .QN(n562) );
  DFFX1 \img_buff_reg[49][3]  ( .D(n4492), .CK(clk), .Q(\img_buff[49][3] ), 
        .QN(n594) );
  DFFX1 \img_buff_reg[53][3]  ( .D(n4524), .CK(clk), .Q(\img_buff[53][3] ), 
        .QN(n626) );
  DFFX1 \img_buff_reg[57][3]  ( .D(n4556), .CK(clk), .Q(\img_buff[57][3] ), 
        .QN(n658) );
  DFFX1 \img_buff_reg[61][3]  ( .D(n4588), .CK(clk), .Q(\img_buff[61][3] ), 
        .QN(n690) );
  DFFX1 \img_buff_reg[3][6]  ( .D(n4121), .CK(clk), .Q(\img_buff[3][6] ), .QN(
        n223) );
  DFFX1 \img_buff_reg[7][6]  ( .D(n4153), .CK(clk), .Q(\img_buff[7][6] ), .QN(
        n255) );
  DFFX1 \img_buff_reg[11][6]  ( .D(n4185), .CK(clk), .Q(\img_buff[11][6] ), 
        .QN(n287) );
  DFFX1 \img_buff_reg[15][6]  ( .D(n4217), .CK(clk), .Q(\img_buff[15][6] ), 
        .QN(n319) );
  DFFX1 \img_buff_reg[19][6]  ( .D(n4249), .CK(clk), .Q(\img_buff[19][6] ), 
        .QN(n351) );
  DFFX1 \img_buff_reg[23][6]  ( .D(n4281), .CK(clk), .Q(\img_buff[23][6] ), 
        .QN(n383) );
  DFFX1 \img_buff_reg[27][6]  ( .D(n4313), .CK(clk), .Q(\img_buff[27][6] ), 
        .QN(n415) );
  DFFX1 \img_buff_reg[31][6]  ( .D(n4345), .CK(clk), .Q(\img_buff[31][6] ), 
        .QN(n447) );
  DFFX1 \img_buff_reg[35][6]  ( .D(n4377), .CK(clk), .Q(\img_buff[35][6] ), 
        .QN(n479) );
  DFFX1 \img_buff_reg[39][6]  ( .D(n4409), .CK(clk), .Q(\img_buff[39][6] ), 
        .QN(n511) );
  DFFX1 \img_buff_reg[43][6]  ( .D(n4441), .CK(clk), .Q(\img_buff[43][6] ), 
        .QN(n543) );
  DFFX1 \img_buff_reg[47][6]  ( .D(n4473), .CK(clk), .Q(\img_buff[47][6] ), 
        .QN(n575) );
  DFFX1 \img_buff_reg[51][6]  ( .D(n4505), .CK(clk), .Q(\img_buff[51][6] ), 
        .QN(n607) );
  DFFX1 \img_buff_reg[55][6]  ( .D(n4537), .CK(clk), .Q(\img_buff[55][6] ), 
        .QN(n639) );
  DFFX1 \img_buff_reg[59][6]  ( .D(n4569), .CK(clk), .Q(\img_buff[59][6] ), 
        .QN(n671) );
  DFFX1 \img_buff_reg[63][6]  ( .D(n4601), .CK(clk), .Q(\img_buff[63][6] ), 
        .QN(n703) );
  DFFX1 \img_buff_reg[7][7]  ( .D(n4152), .CK(clk), .Q(\img_buff[7][7] ), .QN(
        n254) );
  DFFX1 \img_buff_reg[15][7]  ( .D(n4216), .CK(clk), .Q(\img_buff[15][7] ), 
        .QN(n318) );
  DFFX1 \img_buff_reg[19][7]  ( .D(n4248), .CK(clk), .Q(\img_buff[19][7] ), 
        .QN(n350) );
  DFFX1 \img_buff_reg[23][7]  ( .D(n4280), .CK(clk), .Q(\img_buff[23][7] ), 
        .QN(n382) );
  DFFX1 \img_buff_reg[27][7]  ( .D(n4312), .CK(clk), .Q(\img_buff[27][7] ), 
        .QN(n414) );
  DFFX1 \img_buff_reg[31][7]  ( .D(n4344), .CK(clk), .Q(\img_buff[31][7] ), 
        .QN(n446) );
  DFFX1 \img_buff_reg[39][7]  ( .D(n4408), .CK(clk), .Q(\img_buff[39][7] ), 
        .QN(n510) );
  DFFX1 \img_buff_reg[47][7]  ( .D(n4472), .CK(clk), .Q(\img_buff[47][7] ), 
        .QN(n574) );
  DFFX1 \img_buff_reg[51][7]  ( .D(n4504), .CK(clk), .Q(\img_buff[51][7] ), 
        .QN(n606) );
  DFFX1 \img_buff_reg[55][7]  ( .D(n4536), .CK(clk), .Q(\img_buff[55][7] ), 
        .QN(n638) );
  DFFX1 \img_buff_reg[59][7]  ( .D(n4568), .CK(clk), .Q(\img_buff[59][7] ), 
        .QN(n670) );
  DFFX1 \img_buff_reg[63][7]  ( .D(n4600), .CK(clk), .Q(\img_buff[63][7] ), 
        .QN(n702) );
  DFFX1 \img_buff_reg[3][5]  ( .D(n4122), .CK(clk), .Q(\img_buff[3][5] ), .QN(
        n224) );
  DFFX1 \img_buff_reg[7][5]  ( .D(n4154), .CK(clk), .Q(\img_buff[7][5] ), .QN(
        n256) );
  DFFX1 \img_buff_reg[11][5]  ( .D(n4186), .CK(clk), .Q(\img_buff[11][5] ), 
        .QN(n288) );
  DFFX1 \img_buff_reg[15][5]  ( .D(n4218), .CK(clk), .Q(\img_buff[15][5] ), 
        .QN(n320) );
  DFFX1 \img_buff_reg[19][5]  ( .D(n4250), .CK(clk), .Q(\img_buff[19][5] ), 
        .QN(n352) );
  DFFX1 \img_buff_reg[23][5]  ( .D(n4282), .CK(clk), .Q(\img_buff[23][5] ), 
        .QN(n384) );
  DFFX1 \img_buff_reg[27][5]  ( .D(n4314), .CK(clk), .Q(\img_buff[27][5] ), 
        .QN(n416) );
  DFFX1 \img_buff_reg[31][5]  ( .D(n4346), .CK(clk), .Q(\img_buff[31][5] ), 
        .QN(n448) );
  DFFX1 \img_buff_reg[35][5]  ( .D(n4378), .CK(clk), .Q(\img_buff[35][5] ), 
        .QN(n480) );
  DFFX1 \img_buff_reg[39][5]  ( .D(n4410), .CK(clk), .Q(\img_buff[39][5] ), 
        .QN(n512) );
  DFFX1 \img_buff_reg[43][5]  ( .D(n4442), .CK(clk), .Q(\img_buff[43][5] ), 
        .QN(n544) );
  DFFX1 \img_buff_reg[47][5]  ( .D(n4474), .CK(clk), .Q(\img_buff[47][5] ), 
        .QN(n576) );
  DFFX1 \img_buff_reg[51][5]  ( .D(n4506), .CK(clk), .Q(\img_buff[51][5] ), 
        .QN(n608) );
  DFFX1 \img_buff_reg[55][5]  ( .D(n4538), .CK(clk), .Q(\img_buff[55][5] ), 
        .QN(n640) );
  DFFX1 \img_buff_reg[59][5]  ( .D(n4570), .CK(clk), .Q(\img_buff[59][5] ), 
        .QN(n672) );
  DFFX1 \img_buff_reg[63][5]  ( .D(n4602), .CK(clk), .Q(\img_buff[63][5] ), 
        .QN(n704) );
  DFFX1 \img_buff_reg[3][3]  ( .D(n4124), .CK(clk), .Q(\img_buff[3][3] ), .QN(
        n226) );
  DFFX1 \img_buff_reg[7][3]  ( .D(n4156), .CK(clk), .Q(\img_buff[7][3] ), .QN(
        n258) );
  DFFX1 \img_buff_reg[11][3]  ( .D(n4188), .CK(clk), .Q(\img_buff[11][3] ), 
        .QN(n290) );
  DFFX1 \img_buff_reg[15][3]  ( .D(n4220), .CK(clk), .Q(\img_buff[15][3] ), 
        .QN(n322) );
  DFFX1 \img_buff_reg[19][3]  ( .D(n4252), .CK(clk), .Q(\img_buff[19][3] ), 
        .QN(n354) );
  DFFX1 \img_buff_reg[23][3]  ( .D(n4284), .CK(clk), .Q(\img_buff[23][3] ), 
        .QN(n386) );
  DFFX1 \img_buff_reg[27][3]  ( .D(n4316), .CK(clk), .Q(\img_buff[27][3] ), 
        .QN(n418) );
  DFFX1 \img_buff_reg[31][3]  ( .D(n4348), .CK(clk), .Q(\img_buff[31][3] ), 
        .QN(n450) );
  DFFX1 \img_buff_reg[35][3]  ( .D(n4380), .CK(clk), .Q(\img_buff[35][3] ), 
        .QN(n482) );
  DFFX1 \img_buff_reg[39][3]  ( .D(n4412), .CK(clk), .Q(\img_buff[39][3] ), 
        .QN(n514) );
  DFFX1 \img_buff_reg[43][3]  ( .D(n4444), .CK(clk), .Q(\img_buff[43][3] ), 
        .QN(n546) );
  DFFX1 \img_buff_reg[47][3]  ( .D(n4476), .CK(clk), .Q(\img_buff[47][3] ), 
        .QN(n578) );
  DFFX1 \img_buff_reg[51][3]  ( .D(n4508), .CK(clk), .Q(\img_buff[51][3] ), 
        .QN(n610) );
  DFFX1 \img_buff_reg[55][3]  ( .D(n4540), .CK(clk), .Q(\img_buff[55][3] ), 
        .QN(n642) );
  DFFX1 \img_buff_reg[59][3]  ( .D(n4572), .CK(clk), .Q(\img_buff[59][3] ), 
        .QN(n674) );
  DFFX1 \img_buff_reg[63][3]  ( .D(n4604), .CK(clk), .Q(\img_buff[63][3] ), 
        .QN(n706) );
  DFFX1 \img_buff_reg[4][6]  ( .D(n4129), .CK(clk), .Q(\img_buff[4][6] ), .QN(
        n231) );
  DFFX1 \img_buff_reg[8][6]  ( .D(n4161), .CK(clk), .Q(\img_buff[8][6] ), .QN(
        n263) );
  DFFX1 \img_buff_reg[12][6]  ( .D(n4193), .CK(clk), .Q(\img_buff[12][6] ), 
        .QN(n295) );
  DFFX1 \img_buff_reg[16][6]  ( .D(n4225), .CK(clk), .Q(\img_buff[16][6] ), 
        .QN(n327) );
  DFFX1 \img_buff_reg[20][6]  ( .D(n4257), .CK(clk), .Q(\img_buff[20][6] ), 
        .QN(n359) );
  DFFX1 \img_buff_reg[24][6]  ( .D(n4289), .CK(clk), .Q(\img_buff[24][6] ), 
        .QN(n391) );
  DFFX1 \img_buff_reg[28][6]  ( .D(n4321), .CK(clk), .Q(\img_buff[28][6] ), 
        .QN(n423) );
  DFFX1 \img_buff_reg[32][6]  ( .D(n4353), .CK(clk), .Q(\img_buff[32][6] ), 
        .QN(n455) );
  DFFX1 \img_buff_reg[36][6]  ( .D(n4385), .CK(clk), .Q(\img_buff[36][6] ), 
        .QN(n487) );
  DFFX1 \img_buff_reg[40][6]  ( .D(n4417), .CK(clk), .Q(\img_buff[40][6] ), 
        .QN(n519) );
  DFFX1 \img_buff_reg[44][6]  ( .D(n4449), .CK(clk), .Q(\img_buff[44][6] ), 
        .QN(n551) );
  DFFX1 \img_buff_reg[48][6]  ( .D(n4481), .CK(clk), .Q(\img_buff[48][6] ), 
        .QN(n583) );
  DFFX1 \img_buff_reg[52][6]  ( .D(n4513), .CK(clk), .Q(\img_buff[52][6] ), 
        .QN(n615) );
  DFFX1 \img_buff_reg[56][6]  ( .D(n4545), .CK(clk), .Q(\img_buff[56][6] ), 
        .QN(n647) );
  DFFX1 \img_buff_reg[60][6]  ( .D(n4577), .CK(clk), .Q(\img_buff[60][6] ), 
        .QN(n679) );
  DFFX1 \img_buff_reg[20][7]  ( .D(n4256), .CK(clk), .Q(\img_buff[20][7] ), 
        .QN(n358) );
  DFFX1 \img_buff_reg[28][7]  ( .D(n4320), .CK(clk), .Q(\img_buff[28][7] ), 
        .QN(n422) );
  DFFX1 \img_buff_reg[52][7]  ( .D(n4512), .CK(clk), .Q(\img_buff[52][7] ), 
        .QN(n614) );
  DFFX1 \img_buff_reg[60][7]  ( .D(n4576), .CK(clk), .Q(\img_buff[60][7] ), 
        .QN(n678) );
  DFFX1 \img_buff_reg[4][5]  ( .D(n4130), .CK(clk), .Q(\img_buff[4][5] ), .QN(
        n232) );
  DFFX1 \img_buff_reg[8][5]  ( .D(n4162), .CK(clk), .Q(\img_buff[8][5] ), .QN(
        n264) );
  DFFX1 \img_buff_reg[12][5]  ( .D(n4194), .CK(clk), .Q(\img_buff[12][5] ), 
        .QN(n296) );
  DFFX1 \img_buff_reg[16][5]  ( .D(n4226), .CK(clk), .Q(\img_buff[16][5] ), 
        .QN(n328) );
  DFFX1 \img_buff_reg[20][5]  ( .D(n4258), .CK(clk), .Q(\img_buff[20][5] ), 
        .QN(n360) );
  DFFX1 \img_buff_reg[24][5]  ( .D(n4290), .CK(clk), .Q(\img_buff[24][5] ), 
        .QN(n392) );
  DFFX1 \img_buff_reg[28][5]  ( .D(n4322), .CK(clk), .Q(\img_buff[28][5] ), 
        .QN(n424) );
  DFFX1 \img_buff_reg[32][5]  ( .D(n4354), .CK(clk), .Q(\img_buff[32][5] ), 
        .QN(n456) );
  DFFX1 \img_buff_reg[36][5]  ( .D(n4386), .CK(clk), .Q(\img_buff[36][5] ), 
        .QN(n488) );
  DFFX1 \img_buff_reg[40][5]  ( .D(n4418), .CK(clk), .Q(\img_buff[40][5] ), 
        .QN(n520) );
  DFFX1 \img_buff_reg[44][5]  ( .D(n4450), .CK(clk), .Q(\img_buff[44][5] ), 
        .QN(n552) );
  DFFX1 \img_buff_reg[48][5]  ( .D(n4482), .CK(clk), .Q(\img_buff[48][5] ), 
        .QN(n584) );
  DFFX1 \img_buff_reg[52][5]  ( .D(n4514), .CK(clk), .Q(\img_buff[52][5] ), 
        .QN(n616) );
  DFFX1 \img_buff_reg[56][5]  ( .D(n4546), .CK(clk), .Q(\img_buff[56][5] ), 
        .QN(n648) );
  DFFX1 \img_buff_reg[60][5]  ( .D(n4578), .CK(clk), .Q(\img_buff[60][5] ), 
        .QN(n680) );
  DFFX1 \img_buff_reg[4][3]  ( .D(n4132), .CK(clk), .Q(\img_buff[4][3] ), .QN(
        n234) );
  DFFX1 \img_buff_reg[8][3]  ( .D(n4164), .CK(clk), .Q(\img_buff[8][3] ), .QN(
        n266) );
  DFFX1 \img_buff_reg[12][3]  ( .D(n4196), .CK(clk), .Q(\img_buff[12][3] ), 
        .QN(n298) );
  DFFX1 \img_buff_reg[16][3]  ( .D(n4228), .CK(clk), .Q(\img_buff[16][3] ), 
        .QN(n330) );
  DFFX1 \img_buff_reg[20][3]  ( .D(n4260), .CK(clk), .Q(\img_buff[20][3] ), 
        .QN(n362) );
  DFFX1 \img_buff_reg[24][3]  ( .D(n4292), .CK(clk), .Q(\img_buff[24][3] ), 
        .QN(n394) );
  DFFX1 \img_buff_reg[28][3]  ( .D(n4324), .CK(clk), .Q(\img_buff[28][3] ), 
        .QN(n426) );
  DFFX1 \img_buff_reg[32][3]  ( .D(n4356), .CK(clk), .Q(\img_buff[32][3] ), 
        .QN(n458) );
  DFFX1 \img_buff_reg[36][3]  ( .D(n4388), .CK(clk), .Q(\img_buff[36][3] ), 
        .QN(n490) );
  DFFX1 \img_buff_reg[40][3]  ( .D(n4420), .CK(clk), .Q(\img_buff[40][3] ), 
        .QN(n522) );
  DFFX1 \img_buff_reg[44][3]  ( .D(n4452), .CK(clk), .Q(\img_buff[44][3] ), 
        .QN(n554) );
  DFFX1 \img_buff_reg[48][3]  ( .D(n4484), .CK(clk), .Q(\img_buff[48][3] ), 
        .QN(n586) );
  DFFX1 \img_buff_reg[52][3]  ( .D(n4516), .CK(clk), .Q(\img_buff[52][3] ), 
        .QN(n618) );
  DFFX1 \img_buff_reg[56][3]  ( .D(n4548), .CK(clk), .Q(\img_buff[56][3] ), 
        .QN(n650) );
  DFFX1 \img_buff_reg[60][3]  ( .D(n4580), .CK(clk), .Q(\img_buff[60][3] ), 
        .QN(n682) );
  DFFX1 \img_buff_reg[2][6]  ( .D(n4113), .CK(clk), .Q(\img_buff[2][6] ), .QN(
        n215) );
  DFFX1 \img_buff_reg[6][6]  ( .D(n4145), .CK(clk), .Q(\img_buff[6][6] ), .QN(
        n247) );
  DFFX1 \img_buff_reg[10][6]  ( .D(n4177), .CK(clk), .Q(\img_buff[10][6] ), 
        .QN(n279) );
  DFFX1 \img_buff_reg[14][6]  ( .D(n4209), .CK(clk), .Q(\img_buff[14][6] ), 
        .QN(n311) );
  DFFX1 \img_buff_reg[18][6]  ( .D(n4241), .CK(clk), .Q(\img_buff[18][6] ), 
        .QN(n343) );
  DFFX1 \img_buff_reg[22][6]  ( .D(n4273), .CK(clk), .Q(\img_buff[22][6] ), 
        .QN(n375) );
  DFFX1 \img_buff_reg[26][6]  ( .D(n4305), .CK(clk), .Q(\img_buff[26][6] ), 
        .QN(n407) );
  DFFX1 \img_buff_reg[30][6]  ( .D(n4337), .CK(clk), .Q(\img_buff[30][6] ), 
        .QN(n439) );
  DFFX1 \img_buff_reg[34][6]  ( .D(n4369), .CK(clk), .Q(\img_buff[34][6] ), 
        .QN(n471) );
  DFFX1 \img_buff_reg[38][6]  ( .D(n4401), .CK(clk), .Q(\img_buff[38][6] ), 
        .QN(n503) );
  DFFX1 \img_buff_reg[42][6]  ( .D(n4433), .CK(clk), .Q(\img_buff[42][6] ), 
        .QN(n535) );
  DFFX1 \img_buff_reg[46][6]  ( .D(n4465), .CK(clk), .Q(\img_buff[46][6] ), 
        .QN(n567) );
  DFFX1 \img_buff_reg[50][6]  ( .D(n4497), .CK(clk), .Q(\img_buff[50][6] ), 
        .QN(n599) );
  DFFX1 \img_buff_reg[54][6]  ( .D(n4529), .CK(clk), .Q(\img_buff[54][6] ), 
        .QN(n631) );
  DFFX1 \img_buff_reg[58][6]  ( .D(n4561), .CK(clk), .Q(\img_buff[58][6] ), 
        .QN(n663) );
  DFFX1 \img_buff_reg[62][6]  ( .D(n4593), .CK(clk), .Q(\img_buff[62][6] ), 
        .QN(n695) );
  DFFX1 \img_buff_reg[6][7]  ( .D(n4144), .CK(clk), .Q(\img_buff[6][7] ), .QN(
        n246) );
  DFFX1 \img_buff_reg[14][7]  ( .D(n4208), .CK(clk), .Q(\img_buff[14][7] ), 
        .QN(n310) );
  DFFX1 \img_buff_reg[18][7]  ( .D(n4240), .CK(clk), .Q(\img_buff[18][7] ), 
        .QN(n342) );
  DFFX1 \img_buff_reg[22][7]  ( .D(n4272), .CK(clk), .Q(\img_buff[22][7] ), 
        .QN(n374) );
  DFFX1 \img_buff_reg[26][7]  ( .D(n4304), .CK(clk), .Q(\img_buff[26][7] ), 
        .QN(n406) );
  DFFX1 \img_buff_reg[30][7]  ( .D(n4336), .CK(clk), .Q(\img_buff[30][7] ), 
        .QN(n438) );
  DFFX1 \img_buff_reg[38][7]  ( .D(n4400), .CK(clk), .Q(\img_buff[38][7] ), 
        .QN(n502) );
  DFFX1 \img_buff_reg[46][7]  ( .D(n4464), .CK(clk), .Q(\img_buff[46][7] ), 
        .QN(n566) );
  DFFX1 \img_buff_reg[50][7]  ( .D(n4496), .CK(clk), .Q(\img_buff[50][7] ), 
        .QN(n598) );
  DFFX1 \img_buff_reg[54][7]  ( .D(n4528), .CK(clk), .Q(\img_buff[54][7] ), 
        .QN(n630) );
  DFFX1 \img_buff_reg[58][7]  ( .D(n4560), .CK(clk), .Q(\img_buff[58][7] ), 
        .QN(n662) );
  DFFX1 \img_buff_reg[62][7]  ( .D(n4592), .CK(clk), .Q(\img_buff[62][7] ), 
        .QN(n694) );
  DFFX1 \img_buff_reg[2][5]  ( .D(n4114), .CK(clk), .Q(\img_buff[2][5] ), .QN(
        n216) );
  DFFX1 \img_buff_reg[6][5]  ( .D(n4146), .CK(clk), .Q(\img_buff[6][5] ), .QN(
        n248) );
  DFFX1 \img_buff_reg[10][5]  ( .D(n4178), .CK(clk), .Q(\img_buff[10][5] ), 
        .QN(n280) );
  DFFX1 \img_buff_reg[14][5]  ( .D(n4210), .CK(clk), .Q(\img_buff[14][5] ), 
        .QN(n312) );
  DFFX1 \img_buff_reg[18][5]  ( .D(n4242), .CK(clk), .Q(\img_buff[18][5] ), 
        .QN(n344) );
  DFFX1 \img_buff_reg[22][5]  ( .D(n4274), .CK(clk), .Q(\img_buff[22][5] ), 
        .QN(n376) );
  DFFX1 \img_buff_reg[26][5]  ( .D(n4306), .CK(clk), .Q(\img_buff[26][5] ), 
        .QN(n408) );
  DFFX1 \img_buff_reg[30][5]  ( .D(n4338), .CK(clk), .Q(\img_buff[30][5] ), 
        .QN(n440) );
  DFFX1 \img_buff_reg[34][5]  ( .D(n4370), .CK(clk), .Q(\img_buff[34][5] ), 
        .QN(n472) );
  DFFX1 \img_buff_reg[38][5]  ( .D(n4402), .CK(clk), .Q(\img_buff[38][5] ), 
        .QN(n504) );
  DFFX1 \img_buff_reg[42][5]  ( .D(n4434), .CK(clk), .Q(\img_buff[42][5] ), 
        .QN(n536) );
  DFFX1 \img_buff_reg[46][5]  ( .D(n4466), .CK(clk), .Q(\img_buff[46][5] ), 
        .QN(n568) );
  DFFX1 \img_buff_reg[50][5]  ( .D(n4498), .CK(clk), .Q(\img_buff[50][5] ), 
        .QN(n600) );
  DFFX1 \img_buff_reg[54][5]  ( .D(n4530), .CK(clk), .Q(\img_buff[54][5] ), 
        .QN(n632) );
  DFFX1 \img_buff_reg[58][5]  ( .D(n4562), .CK(clk), .Q(\img_buff[58][5] ), 
        .QN(n664) );
  DFFX1 \img_buff_reg[62][5]  ( .D(n4594), .CK(clk), .Q(\img_buff[62][5] ), 
        .QN(n696) );
  DFFX1 \img_buff_reg[2][3]  ( .D(n4116), .CK(clk), .Q(\img_buff[2][3] ), .QN(
        n218) );
  DFFX1 \img_buff_reg[6][3]  ( .D(n4148), .CK(clk), .Q(\img_buff[6][3] ), .QN(
        n250) );
  DFFX1 \img_buff_reg[10][3]  ( .D(n4180), .CK(clk), .Q(\img_buff[10][3] ), 
        .QN(n282) );
  DFFX1 \img_buff_reg[14][3]  ( .D(n4212), .CK(clk), .Q(\img_buff[14][3] ), 
        .QN(n314) );
  DFFX1 \img_buff_reg[18][3]  ( .D(n4244), .CK(clk), .Q(\img_buff[18][3] ), 
        .QN(n346) );
  DFFX1 \img_buff_reg[22][3]  ( .D(n4276), .CK(clk), .Q(\img_buff[22][3] ), 
        .QN(n378) );
  DFFX1 \img_buff_reg[26][3]  ( .D(n4308), .CK(clk), .Q(\img_buff[26][3] ), 
        .QN(n410) );
  DFFX1 \img_buff_reg[30][3]  ( .D(n4340), .CK(clk), .Q(\img_buff[30][3] ), 
        .QN(n442) );
  DFFX1 \img_buff_reg[34][3]  ( .D(n4372), .CK(clk), .Q(\img_buff[34][3] ), 
        .QN(n474) );
  DFFX1 \img_buff_reg[38][3]  ( .D(n4404), .CK(clk), .Q(\img_buff[38][3] ), 
        .QN(n506) );
  DFFX1 \img_buff_reg[42][3]  ( .D(n4436), .CK(clk), .Q(\img_buff[42][3] ), 
        .QN(n538) );
  DFFX1 \img_buff_reg[46][3]  ( .D(n4468), .CK(clk), .Q(\img_buff[46][3] ), 
        .QN(n570) );
  DFFX1 \img_buff_reg[50][3]  ( .D(n4500), .CK(clk), .Q(\img_buff[50][3] ), 
        .QN(n602) );
  DFFX1 \img_buff_reg[54][3]  ( .D(n4532), .CK(clk), .Q(\img_buff[54][3] ), 
        .QN(n634) );
  DFFX1 \img_buff_reg[58][3]  ( .D(n4564), .CK(clk), .Q(\img_buff[58][3] ), 
        .QN(n666) );
  DFFX1 \img_buff_reg[62][3]  ( .D(n4596), .CK(clk), .Q(\img_buff[62][3] ), 
        .QN(n698) );
  DFFQX1 \img_buff_reg[0][7]  ( .D(n6408), .CK(clk), .Q(\img_buff[0][7] ) );
  DFFQX1 \img_buff_reg[0][5]  ( .D(n6409), .CK(clk), .Q(\img_buff[0][5] ) );
  DFFQX1 \img_buff_reg[0][3]  ( .D(n6411), .CK(clk), .Q(\img_buff[0][3] ) );
  DFFX1 \img_buff_reg[1][4]  ( .D(n4107), .CK(clk), .Q(\img_buff[1][4] ), .QN(
        n209) );
  DFFX1 \img_buff_reg[5][4]  ( .D(n4139), .CK(clk), .Q(\img_buff[5][4] ), .QN(
        n241) );
  DFFX1 \img_buff_reg[9][4]  ( .D(n4171), .CK(clk), .Q(\img_buff[9][4] ), .QN(
        n273) );
  DFFX1 \img_buff_reg[13][4]  ( .D(n4203), .CK(clk), .Q(\img_buff[13][4] ), 
        .QN(n305) );
  DFFX1 \img_buff_reg[17][4]  ( .D(n4235), .CK(clk), .Q(\img_buff[17][4] ), 
        .QN(n337) );
  DFFX1 \img_buff_reg[21][4]  ( .D(n4267), .CK(clk), .Q(\img_buff[21][4] ), 
        .QN(n369) );
  DFFX1 \img_buff_reg[25][4]  ( .D(n4299), .CK(clk), .Q(\img_buff[25][4] ), 
        .QN(n401) );
  DFFX1 \img_buff_reg[29][4]  ( .D(n4331), .CK(clk), .Q(\img_buff[29][4] ), 
        .QN(n433) );
  DFFX1 \img_buff_reg[33][4]  ( .D(n4363), .CK(clk), .Q(\img_buff[33][4] ), 
        .QN(n465) );
  DFFX1 \img_buff_reg[37][4]  ( .D(n4395), .CK(clk), .Q(\img_buff[37][4] ), 
        .QN(n497) );
  DFFX1 \img_buff_reg[41][4]  ( .D(n4427), .CK(clk), .Q(\img_buff[41][4] ), 
        .QN(n529) );
  DFFX1 \img_buff_reg[45][4]  ( .D(n4459), .CK(clk), .Q(\img_buff[45][4] ), 
        .QN(n561) );
  DFFX1 \img_buff_reg[49][4]  ( .D(n4491), .CK(clk), .Q(\img_buff[49][4] ), 
        .QN(n593) );
  DFFX1 \img_buff_reg[53][4]  ( .D(n4523), .CK(clk), .Q(\img_buff[53][4] ), 
        .QN(n625) );
  DFFX1 \img_buff_reg[57][4]  ( .D(n4555), .CK(clk), .Q(\img_buff[57][4] ), 
        .QN(n657) );
  DFFX1 \img_buff_reg[61][4]  ( .D(n4587), .CK(clk), .Q(\img_buff[61][4] ), 
        .QN(n689) );
  DFFX1 \img_buff_reg[1][2]  ( .D(n4109), .CK(clk), .Q(\img_buff[1][2] ), .QN(
        n211) );
  DFFX1 \img_buff_reg[5][2]  ( .D(n4141), .CK(clk), .Q(\img_buff[5][2] ), .QN(
        n243) );
  DFFX1 \img_buff_reg[9][2]  ( .D(n4173), .CK(clk), .Q(\img_buff[9][2] ), .QN(
        n275) );
  DFFX1 \img_buff_reg[13][2]  ( .D(n4205), .CK(clk), .Q(\img_buff[13][2] ), 
        .QN(n307) );
  DFFX1 \img_buff_reg[17][2]  ( .D(n4237), .CK(clk), .Q(\img_buff[17][2] ), 
        .QN(n339) );
  DFFX1 \img_buff_reg[21][2]  ( .D(n4269), .CK(clk), .Q(\img_buff[21][2] ), 
        .QN(n371) );
  DFFX1 \img_buff_reg[25][2]  ( .D(n4301), .CK(clk), .Q(\img_buff[25][2] ), 
        .QN(n403) );
  DFFX1 \img_buff_reg[29][2]  ( .D(n4333), .CK(clk), .Q(\img_buff[29][2] ), 
        .QN(n435) );
  DFFX1 \img_buff_reg[33][2]  ( .D(n4365), .CK(clk), .Q(\img_buff[33][2] ), 
        .QN(n467) );
  DFFX1 \img_buff_reg[37][2]  ( .D(n4397), .CK(clk), .Q(\img_buff[37][2] ), 
        .QN(n499) );
  DFFX1 \img_buff_reg[41][2]  ( .D(n4429), .CK(clk), .Q(\img_buff[41][2] ), 
        .QN(n531) );
  DFFX1 \img_buff_reg[45][2]  ( .D(n4461), .CK(clk), .Q(\img_buff[45][2] ), 
        .QN(n563) );
  DFFX1 \img_buff_reg[49][2]  ( .D(n4493), .CK(clk), .Q(\img_buff[49][2] ), 
        .QN(n595) );
  DFFX1 \img_buff_reg[53][2]  ( .D(n4525), .CK(clk), .Q(\img_buff[53][2] ), 
        .QN(n627) );
  DFFX1 \img_buff_reg[57][2]  ( .D(n4557), .CK(clk), .Q(\img_buff[57][2] ), 
        .QN(n659) );
  DFFX1 \img_buff_reg[61][2]  ( .D(n4589), .CK(clk), .Q(\img_buff[61][2] ), 
        .QN(n691) );
  DFFX1 \img_buff_reg[1][1]  ( .D(n4110), .CK(clk), .Q(\img_buff[1][1] ), .QN(
        n212) );
  DFFX1 \img_buff_reg[5][1]  ( .D(n4142), .CK(clk), .Q(\img_buff[5][1] ), .QN(
        n244) );
  DFFX1 \img_buff_reg[17][1]  ( .D(n4238), .CK(clk), .Q(\img_buff[17][1] ), 
        .QN(n340) );
  DFFX1 \img_buff_reg[21][1]  ( .D(n4270), .CK(clk), .Q(\img_buff[21][1] ), 
        .QN(n372) );
  DFFX1 \img_buff_reg[25][1]  ( .D(n4302), .CK(clk), .Q(\img_buff[25][1] ), 
        .QN(n404) );
  DFFX1 \img_buff_reg[29][1]  ( .D(n4334), .CK(clk), .Q(\img_buff[29][1] ), 
        .QN(n436) );
  DFFX1 \img_buff_reg[33][1]  ( .D(n4366), .CK(clk), .Q(\img_buff[33][1] ), 
        .QN(n468) );
  DFFX1 \img_buff_reg[37][1]  ( .D(n4398), .CK(clk), .Q(\img_buff[37][1] ), 
        .QN(n500) );
  DFFX1 \img_buff_reg[41][1]  ( .D(n4430), .CK(clk), .Q(\img_buff[41][1] ), 
        .QN(n532) );
  DFFX1 \img_buff_reg[45][1]  ( .D(n4462), .CK(clk), .Q(\img_buff[45][1] ), 
        .QN(n564) );
  DFFX1 \img_buff_reg[49][1]  ( .D(n4494), .CK(clk), .Q(\img_buff[49][1] ), 
        .QN(n596) );
  DFFX1 \img_buff_reg[53][1]  ( .D(n4526), .CK(clk), .Q(\img_buff[53][1] ), 
        .QN(n628) );
  DFFX1 \img_buff_reg[57][1]  ( .D(n4558), .CK(clk), .Q(\img_buff[57][1] ), 
        .QN(n660) );
  DFFX1 \img_buff_reg[61][1]  ( .D(n4590), .CK(clk), .Q(\img_buff[61][1] ), 
        .QN(n692) );
  DFFX1 \img_buff_reg[1][0]  ( .D(n4111), .CK(clk), .Q(\img_buff[1][0] ), .QN(
        n213) );
  DFFX1 \img_buff_reg[5][0]  ( .D(n4143), .CK(clk), .Q(\img_buff[5][0] ), .QN(
        n245) );
  DFFX1 \img_buff_reg[13][0]  ( .D(n4207), .CK(clk), .Q(\img_buff[13][0] ), 
        .QN(n309) );
  DFFX1 \img_buff_reg[17][0]  ( .D(n4239), .CK(clk), .Q(\img_buff[17][0] ), 
        .QN(n341) );
  DFFX1 \img_buff_reg[21][0]  ( .D(n4271), .CK(clk), .Q(\img_buff[21][0] ), 
        .QN(n373) );
  DFFX1 \img_buff_reg[25][0]  ( .D(n4303), .CK(clk), .Q(\img_buff[25][0] ), 
        .QN(n405) );
  DFFX1 \img_buff_reg[29][0]  ( .D(n4335), .CK(clk), .Q(\img_buff[29][0] ), 
        .QN(n437) );
  DFFX1 \img_buff_reg[33][0]  ( .D(n4367), .CK(clk), .Q(\img_buff[33][0] ), 
        .QN(n469) );
  DFFX1 \img_buff_reg[37][0]  ( .D(n4399), .CK(clk), .Q(\img_buff[37][0] ), 
        .QN(n501) );
  DFFX1 \img_buff_reg[41][0]  ( .D(n4431), .CK(clk), .Q(\img_buff[41][0] ), 
        .QN(n533) );
  DFFX1 \img_buff_reg[45][0]  ( .D(n4463), .CK(clk), .Q(\img_buff[45][0] ), 
        .QN(n565) );
  DFFX1 \img_buff_reg[49][0]  ( .D(n4495), .CK(clk), .Q(\img_buff[49][0] ), 
        .QN(n597) );
  DFFX1 \img_buff_reg[53][0]  ( .D(n4527), .CK(clk), .Q(\img_buff[53][0] ), 
        .QN(n629) );
  DFFX1 \img_buff_reg[61][0]  ( .D(n4591), .CK(clk), .Q(\img_buff[61][0] ), 
        .QN(n693) );
  DFFX1 \img_buff_reg[3][4]  ( .D(n4123), .CK(clk), .Q(\img_buff[3][4] ), .QN(
        n225) );
  DFFX1 \img_buff_reg[11][4]  ( .D(n4187), .CK(clk), .Q(\img_buff[11][4] ), 
        .QN(n289) );
  DFFX1 \img_buff_reg[15][4]  ( .D(n4219), .CK(clk), .Q(\img_buff[15][4] ), 
        .QN(n321) );
  DFFX1 \img_buff_reg[19][4]  ( .D(n4251), .CK(clk), .Q(\img_buff[19][4] ), 
        .QN(n353) );
  DFFX1 \img_buff_reg[23][4]  ( .D(n4283), .CK(clk), .Q(\img_buff[23][4] ), 
        .QN(n385) );
  DFFX1 \img_buff_reg[27][4]  ( .D(n4315), .CK(clk), .Q(\img_buff[27][4] ), 
        .QN(n417) );
  DFFX1 \img_buff_reg[31][4]  ( .D(n4347), .CK(clk), .Q(\img_buff[31][4] ), 
        .QN(n449) );
  DFFX1 \img_buff_reg[35][4]  ( .D(n4379), .CK(clk), .Q(\img_buff[35][4] ), 
        .QN(n481) );
  DFFX1 \img_buff_reg[39][4]  ( .D(n4411), .CK(clk), .Q(\img_buff[39][4] ), 
        .QN(n513) );
  DFFX1 \img_buff_reg[43][4]  ( .D(n4443), .CK(clk), .Q(\img_buff[43][4] ), 
        .QN(n545) );
  DFFX1 \img_buff_reg[47][4]  ( .D(n4475), .CK(clk), .Q(\img_buff[47][4] ), 
        .QN(n577) );
  DFFX1 \img_buff_reg[51][4]  ( .D(n4507), .CK(clk), .Q(\img_buff[51][4] ), 
        .QN(n609) );
  DFFX1 \img_buff_reg[55][4]  ( .D(n4539), .CK(clk), .Q(\img_buff[55][4] ), 
        .QN(n641) );
  DFFX1 \img_buff_reg[59][4]  ( .D(n4571), .CK(clk), .Q(\img_buff[59][4] ), 
        .QN(n673) );
  DFFX1 \img_buff_reg[63][4]  ( .D(n4603), .CK(clk), .Q(\img_buff[63][4] ), 
        .QN(n705) );
  DFFX1 \img_buff_reg[3][2]  ( .D(n4125), .CK(clk), .Q(\img_buff[3][2] ), .QN(
        n227) );
  DFFX1 \img_buff_reg[7][2]  ( .D(n4157), .CK(clk), .Q(\img_buff[7][2] ), .QN(
        n259) );
  DFFX1 \img_buff_reg[11][2]  ( .D(n4189), .CK(clk), .Q(\img_buff[11][2] ), 
        .QN(n291) );
  DFFX1 \img_buff_reg[15][2]  ( .D(n4221), .CK(clk), .Q(\img_buff[15][2] ), 
        .QN(n323) );
  DFFX1 \img_buff_reg[19][2]  ( .D(n4253), .CK(clk), .Q(\img_buff[19][2] ), 
        .QN(n355) );
  DFFX1 \img_buff_reg[23][2]  ( .D(n4285), .CK(clk), .Q(\img_buff[23][2] ), 
        .QN(n387) );
  DFFX1 \img_buff_reg[27][2]  ( .D(n4317), .CK(clk), .Q(\img_buff[27][2] ), 
        .QN(n419) );
  DFFX1 \img_buff_reg[31][2]  ( .D(n4349), .CK(clk), .Q(\img_buff[31][2] ), 
        .QN(n451) );
  DFFX1 \img_buff_reg[35][2]  ( .D(n4381), .CK(clk), .Q(\img_buff[35][2] ), 
        .QN(n483) );
  DFFX1 \img_buff_reg[39][2]  ( .D(n4413), .CK(clk), .Q(\img_buff[39][2] ), 
        .QN(n515) );
  DFFX1 \img_buff_reg[43][2]  ( .D(n4445), .CK(clk), .Q(\img_buff[43][2] ), 
        .QN(n547) );
  DFFX1 \img_buff_reg[47][2]  ( .D(n4477), .CK(clk), .Q(\img_buff[47][2] ), 
        .QN(n579) );
  DFFX1 \img_buff_reg[51][2]  ( .D(n4509), .CK(clk), .Q(\img_buff[51][2] ), 
        .QN(n611) );
  DFFX1 \img_buff_reg[55][2]  ( .D(n4541), .CK(clk), .Q(\img_buff[55][2] ), 
        .QN(n643) );
  DFFX1 \img_buff_reg[59][2]  ( .D(n4573), .CK(clk), .Q(\img_buff[59][2] ), 
        .QN(n675) );
  DFFX1 \img_buff_reg[63][2]  ( .D(n4605), .CK(clk), .Q(\img_buff[63][2] ), 
        .QN(n707) );
  DFFX1 \img_buff_reg[3][1]  ( .D(n4126), .CK(clk), .Q(\img_buff[3][1] ), .QN(
        n228) );
  DFFX1 \img_buff_reg[7][1]  ( .D(n4158), .CK(clk), .Q(\img_buff[7][1] ), .QN(
        n260) );
  DFFX1 \img_buff_reg[11][1]  ( .D(n4190), .CK(clk), .Q(\img_buff[11][1] ), 
        .QN(n292) );
  DFFX1 \img_buff_reg[15][1]  ( .D(n4222), .CK(clk), .Q(\img_buff[15][1] ), 
        .QN(n324) );
  DFFX1 \img_buff_reg[19][1]  ( .D(n4254), .CK(clk), .Q(\img_buff[19][1] ), 
        .QN(n356) );
  DFFX1 \img_buff_reg[23][1]  ( .D(n4286), .CK(clk), .Q(\img_buff[23][1] ), 
        .QN(n388) );
  DFFX1 \img_buff_reg[27][1]  ( .D(n4318), .CK(clk), .Q(\img_buff[27][1] ), 
        .QN(n420) );
  DFFX1 \img_buff_reg[31][1]  ( .D(n4350), .CK(clk), .Q(\img_buff[31][1] ), 
        .QN(n452) );
  DFFX1 \img_buff_reg[35][1]  ( .D(n4382), .CK(clk), .Q(\img_buff[35][1] ), 
        .QN(n484) );
  DFFX1 \img_buff_reg[39][1]  ( .D(n4414), .CK(clk), .Q(\img_buff[39][1] ), 
        .QN(n516) );
  DFFX1 \img_buff_reg[43][1]  ( .D(n4446), .CK(clk), .Q(\img_buff[43][1] ), 
        .QN(n548) );
  DFFX1 \img_buff_reg[47][1]  ( .D(n4478), .CK(clk), .Q(\img_buff[47][1] ), 
        .QN(n580) );
  DFFX1 \img_buff_reg[51][1]  ( .D(n4510), .CK(clk), .Q(\img_buff[51][1] ), 
        .QN(n612) );
  DFFX1 \img_buff_reg[55][1]  ( .D(n4542), .CK(clk), .Q(\img_buff[55][1] ), 
        .QN(n644) );
  DFFX1 \img_buff_reg[59][1]  ( .D(n4574), .CK(clk), .Q(\img_buff[59][1] ), 
        .QN(n676) );
  DFFX1 \img_buff_reg[63][1]  ( .D(n4606), .CK(clk), .Q(\img_buff[63][1] ), 
        .QN(n708) );
  DFFX1 \img_buff_reg[3][0]  ( .D(n4127), .CK(clk), .Q(\img_buff[3][0] ), .QN(
        n229) );
  DFFX1 \img_buff_reg[7][0]  ( .D(n4159), .CK(clk), .Q(\img_buff[7][0] ), .QN(
        n261) );
  DFFX1 \img_buff_reg[15][0]  ( .D(n4223), .CK(clk), .Q(\img_buff[15][0] ), 
        .QN(n325) );
  DFFX1 \img_buff_reg[19][0]  ( .D(n4255), .CK(clk), .Q(\img_buff[19][0] ), 
        .QN(n357) );
  DFFX1 \img_buff_reg[23][0]  ( .D(n4287), .CK(clk), .Q(\img_buff[23][0] ), 
        .QN(n389) );
  DFFX1 \img_buff_reg[27][0]  ( .D(n4319), .CK(clk), .Q(\img_buff[27][0] ), 
        .QN(n421) );
  DFFX1 \img_buff_reg[31][0]  ( .D(n4351), .CK(clk), .Q(\img_buff[31][0] ), 
        .QN(n453) );
  DFFX1 \img_buff_reg[35][0]  ( .D(n4383), .CK(clk), .Q(\img_buff[35][0] ), 
        .QN(n485) );
  DFFX1 \img_buff_reg[39][0]  ( .D(n4415), .CK(clk), .Q(\img_buff[39][0] ), 
        .QN(n517) );
  DFFX1 \img_buff_reg[43][0]  ( .D(n4447), .CK(clk), .Q(\img_buff[43][0] ), 
        .QN(n549) );
  DFFX1 \img_buff_reg[47][0]  ( .D(n4479), .CK(clk), .Q(\img_buff[47][0] ), 
        .QN(n581) );
  DFFX1 \img_buff_reg[51][0]  ( .D(n4511), .CK(clk), .Q(\img_buff[51][0] ), 
        .QN(n613) );
  DFFX1 \img_buff_reg[59][0]  ( .D(n4575), .CK(clk), .Q(\img_buff[59][0] ), 
        .QN(n677) );
  DFFX1 \img_buff_reg[4][4]  ( .D(n4131), .CK(clk), .Q(\img_buff[4][4] ), .QN(
        n233) );
  DFFX1 \img_buff_reg[12][4]  ( .D(n4195), .CK(clk), .Q(\img_buff[12][4] ), 
        .QN(n297) );
  DFFX1 \img_buff_reg[16][4]  ( .D(n4227), .CK(clk), .Q(\img_buff[16][4] ), 
        .QN(n329) );
  DFFX1 \img_buff_reg[20][4]  ( .D(n4259), .CK(clk), .Q(\img_buff[20][4] ), 
        .QN(n361) );
  DFFX1 \img_buff_reg[24][4]  ( .D(n4291), .CK(clk), .Q(\img_buff[24][4] ), 
        .QN(n393) );
  DFFX1 \img_buff_reg[28][4]  ( .D(n4323), .CK(clk), .Q(\img_buff[28][4] ), 
        .QN(n425) );
  DFFX1 \img_buff_reg[32][4]  ( .D(n4355), .CK(clk), .Q(\img_buff[32][4] ), 
        .QN(n457) );
  DFFX1 \img_buff_reg[36][4]  ( .D(n4387), .CK(clk), .Q(\img_buff[36][4] ), 
        .QN(n489) );
  DFFX1 \img_buff_reg[40][4]  ( .D(n4419), .CK(clk), .Q(\img_buff[40][4] ), 
        .QN(n521) );
  DFFX1 \img_buff_reg[44][4]  ( .D(n4451), .CK(clk), .Q(\img_buff[44][4] ), 
        .QN(n553) );
  DFFX1 \img_buff_reg[48][4]  ( .D(n4483), .CK(clk), .Q(\img_buff[48][4] ), 
        .QN(n585) );
  DFFX1 \img_buff_reg[52][4]  ( .D(n4515), .CK(clk), .Q(\img_buff[52][4] ), 
        .QN(n617) );
  DFFX1 \img_buff_reg[56][4]  ( .D(n4547), .CK(clk), .Q(\img_buff[56][4] ), 
        .QN(n649) );
  DFFX1 \img_buff_reg[60][4]  ( .D(n4579), .CK(clk), .Q(\img_buff[60][4] ), 
        .QN(n681) );
  DFFX1 \img_buff_reg[4][2]  ( .D(n4133), .CK(clk), .Q(\img_buff[4][2] ), .QN(
        n235) );
  DFFX1 \img_buff_reg[8][2]  ( .D(n4165), .CK(clk), .Q(\img_buff[8][2] ), .QN(
        n267) );
  DFFX1 \img_buff_reg[12][2]  ( .D(n4197), .CK(clk), .Q(\img_buff[12][2] ), 
        .QN(n299) );
  DFFX1 \img_buff_reg[16][2]  ( .D(n4229), .CK(clk), .Q(\img_buff[16][2] ), 
        .QN(n331) );
  DFFX1 \img_buff_reg[20][2]  ( .D(n4261), .CK(clk), .Q(\img_buff[20][2] ), 
        .QN(n363) );
  DFFX1 \img_buff_reg[24][2]  ( .D(n4293), .CK(clk), .Q(\img_buff[24][2] ), 
        .QN(n395) );
  DFFX1 \img_buff_reg[28][2]  ( .D(n4325), .CK(clk), .Q(\img_buff[28][2] ), 
        .QN(n427) );
  DFFX1 \img_buff_reg[32][2]  ( .D(n4357), .CK(clk), .Q(\img_buff[32][2] ), 
        .QN(n459) );
  DFFX1 \img_buff_reg[36][2]  ( .D(n4389), .CK(clk), .Q(\img_buff[36][2] ), 
        .QN(n491) );
  DFFX1 \img_buff_reg[40][2]  ( .D(n4421), .CK(clk), .Q(\img_buff[40][2] ), 
        .QN(n523) );
  DFFX1 \img_buff_reg[44][2]  ( .D(n4453), .CK(clk), .Q(\img_buff[44][2] ), 
        .QN(n555) );
  DFFX1 \img_buff_reg[48][2]  ( .D(n4485), .CK(clk), .Q(\img_buff[48][2] ), 
        .QN(n587) );
  DFFX1 \img_buff_reg[52][2]  ( .D(n4517), .CK(clk), .Q(\img_buff[52][2] ), 
        .QN(n619) );
  DFFX1 \img_buff_reg[56][2]  ( .D(n4549), .CK(clk), .Q(\img_buff[56][2] ), 
        .QN(n651) );
  DFFX1 \img_buff_reg[60][2]  ( .D(n4581), .CK(clk), .Q(\img_buff[60][2] ), 
        .QN(n683) );
  DFFX1 \img_buff_reg[4][1]  ( .D(n4134), .CK(clk), .Q(\img_buff[4][1] ), .QN(
        n236) );
  DFFX1 \img_buff_reg[8][1]  ( .D(n4166), .CK(clk), .Q(\img_buff[8][1] ), .QN(
        n268) );
  DFFX1 \img_buff_reg[12][1]  ( .D(n4198), .CK(clk), .Q(\img_buff[12][1] ), 
        .QN(n300) );
  DFFX1 \img_buff_reg[16][1]  ( .D(n4230), .CK(clk), .Q(\img_buff[16][1] ), 
        .QN(n332) );
  DFFX1 \img_buff_reg[20][1]  ( .D(n4262), .CK(clk), .Q(\img_buff[20][1] ), 
        .QN(n364) );
  DFFX1 \img_buff_reg[24][1]  ( .D(n4294), .CK(clk), .Q(\img_buff[24][1] ), 
        .QN(n396) );
  DFFX1 \img_buff_reg[28][1]  ( .D(n4326), .CK(clk), .Q(\img_buff[28][1] ), 
        .QN(n428) );
  DFFX1 \img_buff_reg[32][1]  ( .D(n4358), .CK(clk), .Q(\img_buff[32][1] ), 
        .QN(n460) );
  DFFX1 \img_buff_reg[36][1]  ( .D(n4390), .CK(clk), .Q(\img_buff[36][1] ), 
        .QN(n492) );
  DFFX1 \img_buff_reg[40][1]  ( .D(n4422), .CK(clk), .Q(\img_buff[40][1] ), 
        .QN(n524) );
  DFFX1 \img_buff_reg[44][1]  ( .D(n4454), .CK(clk), .Q(\img_buff[44][1] ), 
        .QN(n556) );
  DFFX1 \img_buff_reg[48][1]  ( .D(n4486), .CK(clk), .Q(\img_buff[48][1] ), 
        .QN(n588) );
  DFFX1 \img_buff_reg[52][1]  ( .D(n4518), .CK(clk), .Q(\img_buff[52][1] ), 
        .QN(n620) );
  DFFX1 \img_buff_reg[56][1]  ( .D(n4550), .CK(clk), .Q(\img_buff[56][1] ), 
        .QN(n652) );
  DFFX1 \img_buff_reg[60][1]  ( .D(n4582), .CK(clk), .Q(\img_buff[60][1] ), 
        .QN(n684) );
  DFFX1 \img_buff_reg[4][0]  ( .D(n4135), .CK(clk), .Q(\img_buff[4][0] ), .QN(
        n237) );
  DFFX1 \img_buff_reg[8][0]  ( .D(n4167), .CK(clk), .Q(\img_buff[8][0] ), .QN(
        n269) );
  DFFX1 \img_buff_reg[12][0]  ( .D(n4199), .CK(clk), .Q(\img_buff[12][0] ), 
        .QN(n301) );
  DFFX1 \img_buff_reg[16][0]  ( .D(n4231), .CK(clk), .Q(\img_buff[16][0] ), 
        .QN(n333) );
  DFFX1 \img_buff_reg[20][0]  ( .D(n4263), .CK(clk), .Q(\img_buff[20][0] ), 
        .QN(n365) );
  DFFX1 \img_buff_reg[24][0]  ( .D(n4295), .CK(clk), .Q(\img_buff[24][0] ), 
        .QN(n397) );
  DFFX1 \img_buff_reg[28][0]  ( .D(n4327), .CK(clk), .Q(\img_buff[28][0] ), 
        .QN(n429) );
  DFFX1 \img_buff_reg[32][0]  ( .D(n4359), .CK(clk), .Q(\img_buff[32][0] ), 
        .QN(n461) );
  DFFX1 \img_buff_reg[36][0]  ( .D(n4391), .CK(clk), .Q(\img_buff[36][0] ), 
        .QN(n493) );
  DFFX1 \img_buff_reg[40][0]  ( .D(n4423), .CK(clk), .Q(\img_buff[40][0] ), 
        .QN(n525) );
  DFFX1 \img_buff_reg[44][0]  ( .D(n4455), .CK(clk), .Q(\img_buff[44][0] ), 
        .QN(n557) );
  DFFX1 \img_buff_reg[48][0]  ( .D(n4487), .CK(clk), .Q(\img_buff[48][0] ), 
        .QN(n589) );
  DFFX1 \img_buff_reg[52][0]  ( .D(n4519), .CK(clk), .Q(\img_buff[52][0] ), 
        .QN(n621) );
  DFFX1 \img_buff_reg[56][0]  ( .D(n4551), .CK(clk), .Q(\img_buff[56][0] ), 
        .QN(n653) );
  DFFX1 \img_buff_reg[60][0]  ( .D(n4583), .CK(clk), .Q(\img_buff[60][0] ), 
        .QN(n685) );
  DFFX1 \img_buff_reg[2][4]  ( .D(n4115), .CK(clk), .Q(\img_buff[2][4] ), .QN(
        n217) );
  DFFX1 \img_buff_reg[6][4]  ( .D(n4147), .CK(clk), .Q(\img_buff[6][4] ), .QN(
        n249) );
  DFFX1 \img_buff_reg[10][4]  ( .D(n4179), .CK(clk), .Q(\img_buff[10][4] ), 
        .QN(n281) );
  DFFX1 \img_buff_reg[14][4]  ( .D(n4211), .CK(clk), .Q(\img_buff[14][4] ), 
        .QN(n313) );
  DFFX1 \img_buff_reg[18][4]  ( .D(n4243), .CK(clk), .Q(\img_buff[18][4] ), 
        .QN(n345) );
  DFFX1 \img_buff_reg[22][4]  ( .D(n4275), .CK(clk), .Q(\img_buff[22][4] ), 
        .QN(n377) );
  DFFX1 \img_buff_reg[26][4]  ( .D(n4307), .CK(clk), .Q(\img_buff[26][4] ), 
        .QN(n409) );
  DFFX1 \img_buff_reg[30][4]  ( .D(n4339), .CK(clk), .Q(\img_buff[30][4] ), 
        .QN(n441) );
  DFFX1 \img_buff_reg[34][4]  ( .D(n4371), .CK(clk), .Q(\img_buff[34][4] ), 
        .QN(n473) );
  DFFX1 \img_buff_reg[38][4]  ( .D(n4403), .CK(clk), .Q(\img_buff[38][4] ), 
        .QN(n505) );
  DFFX1 \img_buff_reg[42][4]  ( .D(n4435), .CK(clk), .Q(\img_buff[42][4] ), 
        .QN(n537) );
  DFFX1 \img_buff_reg[46][4]  ( .D(n4467), .CK(clk), .Q(\img_buff[46][4] ), 
        .QN(n569) );
  DFFX1 \img_buff_reg[50][4]  ( .D(n4499), .CK(clk), .Q(\img_buff[50][4] ), 
        .QN(n601) );
  DFFX1 \img_buff_reg[54][4]  ( .D(n4531), .CK(clk), .Q(\img_buff[54][4] ), 
        .QN(n633) );
  DFFX1 \img_buff_reg[58][4]  ( .D(n4563), .CK(clk), .Q(\img_buff[58][4] ), 
        .QN(n665) );
  DFFX1 \img_buff_reg[62][4]  ( .D(n4595), .CK(clk), .Q(\img_buff[62][4] ), 
        .QN(n697) );
  DFFX1 \img_buff_reg[2][2]  ( .D(n4117), .CK(clk), .Q(\img_buff[2][2] ), .QN(
        n219) );
  DFFX1 \img_buff_reg[6][2]  ( .D(n4149), .CK(clk), .Q(\img_buff[6][2] ), .QN(
        n251) );
  DFFX1 \img_buff_reg[10][2]  ( .D(n4181), .CK(clk), .Q(\img_buff[10][2] ), 
        .QN(n283) );
  DFFX1 \img_buff_reg[14][2]  ( .D(n4213), .CK(clk), .Q(\img_buff[14][2] ), 
        .QN(n315) );
  DFFX1 \img_buff_reg[18][2]  ( .D(n4245), .CK(clk), .Q(\img_buff[18][2] ), 
        .QN(n347) );
  DFFX1 \img_buff_reg[22][2]  ( .D(n4277), .CK(clk), .Q(\img_buff[22][2] ), 
        .QN(n379) );
  DFFX1 \img_buff_reg[26][2]  ( .D(n4309), .CK(clk), .Q(\img_buff[26][2] ), 
        .QN(n411) );
  DFFX1 \img_buff_reg[30][2]  ( .D(n4341), .CK(clk), .Q(\img_buff[30][2] ), 
        .QN(n443) );
  DFFX1 \img_buff_reg[34][2]  ( .D(n4373), .CK(clk), .Q(\img_buff[34][2] ), 
        .QN(n475) );
  DFFX1 \img_buff_reg[38][2]  ( .D(n4405), .CK(clk), .Q(\img_buff[38][2] ), 
        .QN(n507) );
  DFFX1 \img_buff_reg[42][2]  ( .D(n4437), .CK(clk), .Q(\img_buff[42][2] ), 
        .QN(n539) );
  DFFX1 \img_buff_reg[46][2]  ( .D(n4469), .CK(clk), .Q(\img_buff[46][2] ), 
        .QN(n571) );
  DFFX1 \img_buff_reg[50][2]  ( .D(n4501), .CK(clk), .Q(\img_buff[50][2] ), 
        .QN(n603) );
  DFFX1 \img_buff_reg[54][2]  ( .D(n4533), .CK(clk), .Q(\img_buff[54][2] ), 
        .QN(n635) );
  DFFX1 \img_buff_reg[58][2]  ( .D(n4565), .CK(clk), .Q(\img_buff[58][2] ), 
        .QN(n667) );
  DFFX1 \img_buff_reg[62][2]  ( .D(n4597), .CK(clk), .Q(\img_buff[62][2] ), 
        .QN(n699) );
  DFFX1 \img_buff_reg[2][1]  ( .D(n4118), .CK(clk), .Q(\img_buff[2][1] ), .QN(
        n220) );
  DFFX1 \img_buff_reg[6][1]  ( .D(n4150), .CK(clk), .Q(\img_buff[6][1] ), .QN(
        n252) );
  DFFX1 \img_buff_reg[10][1]  ( .D(n4182), .CK(clk), .Q(\img_buff[10][1] ), 
        .QN(n284) );
  DFFX1 \img_buff_reg[14][1]  ( .D(n4214), .CK(clk), .Q(\img_buff[14][1] ), 
        .QN(n316) );
  DFFX1 \img_buff_reg[18][1]  ( .D(n4246), .CK(clk), .Q(\img_buff[18][1] ), 
        .QN(n348) );
  DFFX1 \img_buff_reg[22][1]  ( .D(n4278), .CK(clk), .Q(\img_buff[22][1] ), 
        .QN(n380) );
  DFFX1 \img_buff_reg[26][1]  ( .D(n4310), .CK(clk), .Q(\img_buff[26][1] ), 
        .QN(n412) );
  DFFX1 \img_buff_reg[30][1]  ( .D(n4342), .CK(clk), .Q(\img_buff[30][1] ), 
        .QN(n444) );
  DFFX1 \img_buff_reg[34][1]  ( .D(n4374), .CK(clk), .Q(\img_buff[34][1] ), 
        .QN(n476) );
  DFFX1 \img_buff_reg[38][1]  ( .D(n4406), .CK(clk), .Q(\img_buff[38][1] ), 
        .QN(n508) );
  DFFX1 \img_buff_reg[42][1]  ( .D(n4438), .CK(clk), .Q(\img_buff[42][1] ), 
        .QN(n540) );
  DFFX1 \img_buff_reg[46][1]  ( .D(n4470), .CK(clk), .Q(\img_buff[46][1] ), 
        .QN(n572) );
  DFFX1 \img_buff_reg[50][1]  ( .D(n4502), .CK(clk), .Q(\img_buff[50][1] ), 
        .QN(n604) );
  DFFX1 \img_buff_reg[54][1]  ( .D(n4534), .CK(clk), .Q(\img_buff[54][1] ), 
        .QN(n636) );
  DFFX1 \img_buff_reg[58][1]  ( .D(n4566), .CK(clk), .Q(\img_buff[58][1] ), 
        .QN(n668) );
  DFFX1 \img_buff_reg[62][1]  ( .D(n4598), .CK(clk), .Q(\img_buff[62][1] ), 
        .QN(n700) );
  DFFX1 \img_buff_reg[2][0]  ( .D(n4119), .CK(clk), .Q(\img_buff[2][0] ), .QN(
        n221) );
  DFFX1 \img_buff_reg[6][0]  ( .D(n4151), .CK(clk), .Q(\img_buff[6][0] ), .QN(
        n253) );
  DFFX1 \img_buff_reg[14][0]  ( .D(n4215), .CK(clk), .Q(\img_buff[14][0] ), 
        .QN(n317) );
  DFFX1 \img_buff_reg[18][0]  ( .D(n4247), .CK(clk), .Q(\img_buff[18][0] ), 
        .QN(n349) );
  DFFX1 \img_buff_reg[22][0]  ( .D(n4279), .CK(clk), .Q(\img_buff[22][0] ), 
        .QN(n381) );
  DFFX1 \img_buff_reg[26][0]  ( .D(n4311), .CK(clk), .Q(\img_buff[26][0] ), 
        .QN(n413) );
  DFFX1 \img_buff_reg[30][0]  ( .D(n4343), .CK(clk), .Q(\img_buff[30][0] ), 
        .QN(n445) );
  DFFX1 \img_buff_reg[34][0]  ( .D(n4375), .CK(clk), .Q(\img_buff[34][0] ), 
        .QN(n477) );
  DFFX1 \img_buff_reg[38][0]  ( .D(n4407), .CK(clk), .Q(\img_buff[38][0] ), 
        .QN(n509) );
  DFFX1 \img_buff_reg[42][0]  ( .D(n4439), .CK(clk), .Q(\img_buff[42][0] ), 
        .QN(n541) );
  DFFX1 \img_buff_reg[46][0]  ( .D(n4471), .CK(clk), .Q(\img_buff[46][0] ), 
        .QN(n573) );
  DFFX1 \img_buff_reg[50][0]  ( .D(n4503), .CK(clk), .Q(\img_buff[50][0] ), 
        .QN(n605) );
  DFFX1 \img_buff_reg[54][0]  ( .D(n4535), .CK(clk), .Q(\img_buff[54][0] ), 
        .QN(n637) );
  DFFX1 \img_buff_reg[58][0]  ( .D(n4567), .CK(clk), .Q(\img_buff[58][0] ), 
        .QN(n669) );
  DFFX1 \img_buff_reg[62][0]  ( .D(n4599), .CK(clk), .Q(\img_buff[62][0] ), 
        .QN(n701) );
  DFFQX1 \img_buff_reg[0][4]  ( .D(n6410), .CK(clk), .Q(\img_buff[0][4] ) );
  DFFQX1 \img_buff_reg[0][2]  ( .D(n6412), .CK(clk), .Q(\img_buff[0][2] ) );
  DFFQX1 \img_buff_reg[0][1]  ( .D(n6413), .CK(clk), .Q(\img_buff[0][1] ) );
  DFFQX1 \img_buff_reg[0][0]  ( .D(n6414), .CK(clk), .Q(\img_buff[0][0] ) );
  ADDHXL \add_118/U1_1_4  ( .A(n6673), .B(\add_118/carry[4] ), .CO(
        \add_118/carry[5] ), .S(N3384) );
  ADDHXL \add_139/U1_1_4  ( .A(IRAM_A[4]), .B(\add_139/carry[4] ), .CO(
        \add_139/carry[5] ), .S(N3454) );
  ADDHXL \add_118/U1_1_3  ( .A(n6674), .B(\add_118/carry[3] ), .CO(
        \add_118/carry[4] ), .S(N3383) );
  ADDHXL \add_118/U1_1_2  ( .A(IROM_A[2]), .B(\add_118/carry[2] ), .CO(
        \add_118/carry[3] ), .S(N3382) );
  ADDHXL \add_139/U1_1_2  ( .A(IRAM_A[2]), .B(\add_139/carry[2] ), .CO(
        \add_139/carry[3] ), .S(N3452) );
  ADDHXL \add_139/U1_1_3  ( .A(IRAM_A[3]), .B(\add_139/carry[3] ), .CO(
        \add_139/carry[4] ), .S(N3453) );
  ADDHXL \add_118/U1_1_1  ( .A(IROM_A[1]), .B(n6677), .CO(\add_118/carry[2] ), 
        .S(N3381) );
  ADDHXL \add_139/U1_1_1  ( .A(IRAM_A[1]), .B(n6692), .CO(\add_139/carry[2] ), 
        .S(N3451) );
  DFFHQX8 \col_reg[0]  ( .D(n4610), .CK(clk), .Q(N3323) );
  DFFQX1 \img_buff_reg[0][6]  ( .D(n4672), .CK(clk), .Q(\img_buff[0][6] ) );
  EDFFXL \avg_reg[7]  ( .D(N6166), .E(N16287), .CK(clk), .QN(n162) );
  EDFFXL \avg_reg[6]  ( .D(N6165), .E(N16287), .CK(clk), .QN(n164) );
  EDFFXL \avg_reg[5]  ( .D(N6164), .E(N16287), .CK(clk), .QN(n166) );
  EDFFXL \avg_reg[4]  ( .D(N6163), .E(N16287), .CK(clk), .QN(n168) );
  DFFX1 \img_buff_reg[13][1]  ( .D(n4206), .CK(clk), .Q(\img_buff[13][1] ), 
        .QN(n308) );
  DFFX1 \img_buff_reg[9][1]  ( .D(n4174), .CK(clk), .Q(\img_buff[9][1] ), .QN(
        n276) );
  DFFX1 \img_buff_reg[8][4]  ( .D(n4163), .CK(clk), .Q(\img_buff[8][4] ), .QN(
        n265) );
  DFFQX1 \row_reg[2]  ( .D(n4613), .CK(clk), .Q(N3340) );
  DFFQX2 \IRAM_A_reg[0]  ( .D(n4625), .CK(clk), .Q(n6692) );
  DFFQX2 \IROM_A_reg[0]  ( .D(n4619), .CK(clk), .Q(n6677) );
  DFFQX1 \IRAM_A_reg[5]  ( .D(n4626), .CK(clk), .Q(n6687) );
  DFFQX1 \IRAM_A_reg[2]  ( .D(n4623), .CK(clk), .Q(n6690) );
  DFFQX1 \IRAM_A_reg[4]  ( .D(n4621), .CK(clk), .Q(n6688) );
  DFFQX1 \IROM_A_reg[3]  ( .D(n4616), .CK(clk), .Q(n6674) );
  DFFQX1 IRAM_valid_reg ( .D(n4608), .CK(clk), .Q(n6678) );
  DFFQX1 \IRAM_D_reg[0]  ( .D(n4103), .CK(clk), .Q(n6686) );
  DFFQX1 \IRAM_D_reg[1]  ( .D(n4102), .CK(clk), .Q(n6685) );
  DFFQX1 \IRAM_D_reg[2]  ( .D(n4101), .CK(clk), .Q(n6684) );
  DFFQX1 \IRAM_D_reg[3]  ( .D(n4100), .CK(clk), .Q(n6683) );
  DFFQX1 \IRAM_D_reg[4]  ( .D(n4099), .CK(clk), .Q(n6682) );
  DFFQX1 \IRAM_D_reg[5]  ( .D(n4098), .CK(clk), .Q(n6681) );
  DFFQX1 \IRAM_D_reg[7]  ( .D(n4096), .CK(clk), .Q(n6679) );
  DFFQX1 \IRAM_D_reg[6]  ( .D(n4097), .CK(clk), .Q(n6680) );
  DFFQX1 IROM_rd_reg ( .D(n4614), .CK(clk), .Q(n6671) );
  DFFQX1 \IRAM_A_reg[3]  ( .D(n4622), .CK(clk), .Q(n6689) );
  DFFQX1 \IRAM_A_reg[1]  ( .D(n4624), .CK(clk), .Q(n6691) );
  DFFQX1 \IROM_A_reg[2]  ( .D(n4617), .CK(clk), .Q(n6675) );
  DFFQX1 \IROM_A_reg[5]  ( .D(n4620), .CK(clk), .Q(n6672) );
  DFFQX1 \IROM_A_reg[1]  ( .D(n4618), .CK(clk), .Q(n6676) );
  DFFQX1 \IROM_A_reg[4]  ( .D(n4615), .CK(clk), .Q(n6673) );
  EDFFX1 \cmd_reg_reg[3]  ( .D(cmd[3]), .E(n4883), .CK(clk), .Q(cmd_reg[3]) );
  EDFFX1 \cmd_reg_reg[2]  ( .D(cmd[2]), .E(n4883), .CK(clk), .Q(cmd_reg[2]) );
  EDFFHQX1 busy_reg ( .D(n967), .E(n968), .CK(clk), .Q(n4729) );
  DFFX1 \img_buff_reg[55][0]  ( .D(n4543), .CK(clk), .Q(\img_buff[55][0] ), 
        .QN(n645) );
  DFFX1 \img_buff_reg[10][0]  ( .D(n4183), .CK(clk), .Q(\img_buff[10][0] ), 
        .QN(n285) );
  DFFX1 \img_buff_reg[57][0]  ( .D(n4559), .CK(clk), .Q(\img_buff[57][0] ), 
        .QN(n661) );
  DFFX1 \img_buff_reg[7][4]  ( .D(n4155), .CK(clk), .Q(\img_buff[7][4] ), .QN(
        n257) );
  DFFX1 \img_buff_reg[9][0]  ( .D(n4175), .CK(clk), .Q(\img_buff[9][0] ), .QN(
        n277) );
  DFFX1 \img_buff_reg[11][0]  ( .D(n4191), .CK(clk), .Q(\img_buff[11][0] ), 
        .QN(n293) );
  DFFX1 \img_buff_reg[63][0]  ( .D(n4607), .CK(clk), .Q(\img_buff[63][0] ), 
        .QN(n709) );
  DFFQX2 \row_reg[1]  ( .D(n4611), .CK(clk), .Q(N3339) );
  DFFQX2 \row_reg[0]  ( .D(n4612), .CK(clk), .Q(N3338) );
  EDFFX2 \col_reg[2]  ( .D(n6643), .E(n4064), .CK(clk), .Q(N3325), .QN(n944)
         );
  DFFHQX4 \col_reg[1]  ( .D(n4609), .CK(clk), .Q(N3324) );
  BUFX2 U4062 ( .A(n5082), .Y(n5072) );
  BUFX12 U4063 ( .A(n1040), .Y(n4627) );
  BUFX4 U4064 ( .A(n5071), .Y(n5075) );
  CLKBUFX2 U4065 ( .A(n5082), .Y(n5071) );
  CLKBUFX3 U4066 ( .A(n5791), .Y(n4628) );
  CLKBUFX3 U4067 ( .A(n5791), .Y(n4629) );
  CLKBUFX3 U4068 ( .A(n5791), .Y(n4630) );
  INVX2 U4069 ( .A(n5796), .Y(n5791) );
  INVX6 U4070 ( .A(n5923), .Y(n5920) );
  CLKBUFX4 U4071 ( .A(n5638), .Y(n5640) );
  BUFX3 U4072 ( .A(n5638), .Y(n5639) );
  CLKBUFX2 U4073 ( .A(n5970), .Y(n4631) );
  CLKBUFX2 U4074 ( .A(n5970), .Y(n4632) );
  CLKINVX1 U4075 ( .A(n4695), .Y(n4633) );
  CLKINVX1 U4076 ( .A(n5055), .Y(n4634) );
  INVXL U4077 ( .A(n5062), .Y(n4635) );
  INVXL U4078 ( .A(n4762), .Y(n4636) );
  CLKBUFX3 U4079 ( .A(n5064), .Y(n5055) );
  BUFX12 U4080 ( .A(n5056), .Y(n5063) );
  XOR2X1 U4081 ( .A(N3324), .B(N3323), .Y(n4805) );
  CLKINVX12 U4082 ( .A(n4762), .Y(n4763) );
  CLKBUFX3 U4083 ( .A(n5254), .Y(n5247) );
  INVX8 U4084 ( .A(n1037), .Y(n5796) );
  OAI222X2 U4085 ( .A0(n3998), .A1(n3975), .B0(n3999), .B1(n5668), .C0(n4000), 
        .C1(n162), .Y(n997) );
  AOI221X1 U4086 ( .A0(n5659), .A1(n3982), .B0(n5941), .B1(n3983), .C0(n4002), 
        .Y(n3998) );
  BUFX16 U4087 ( .A(n1048), .Y(n4637) );
  MX4X1 U4088 ( .A(n4918), .B(n4916), .C(n4917), .D(n4915), .S0(n5067), .S1(
        n5065), .Y(n4919) );
  BUFX6 U4089 ( .A(n5069), .Y(n5067) );
  CLKBUFX8 U4090 ( .A(n5246), .Y(n5250) );
  NOR2BX2 U4091 ( .AN(n5457), .B(n5666), .Y(n6231) );
  OAI31X4 U4092 ( .A0(n6224), .A1(n6223), .A2(n6222), .B0(n6221), .Y(N5342) );
  CLKINVX1 U4093 ( .A(n6046), .Y(n6069) );
  NOR3BX1 U4094 ( .AN(n6060), .B(n6059), .C(n6045), .Y(n6046) );
  OAI2BB1X4 U4095 ( .A0N(n4053), .A1N(n4035), .B0(n4036), .Y(n1053) );
  BUFX12 U4096 ( .A(n1053), .Y(n5785) );
  AOI31X1 U4097 ( .A0(n6090), .A1(n6089), .A2(n6088), .B0(n6087), .Y(n6094) );
  NOR2BX2 U4098 ( .AN(N3359), .B(n5457), .Y(n6291) );
  NOR2BX4 U4099 ( .AN(n5666), .B(n5457), .Y(n6319) );
  MX4X4 U4100 ( .A(n5483), .B(n5473), .C(n5478), .D(n5468), .S0(n5672), .S1(
        n5674), .Y(n5457) );
  BUFX4 U4101 ( .A(n5789), .Y(n4638) );
  BUFX6 U4102 ( .A(n5789), .Y(n4639) );
  CLKBUFX4 U4103 ( .A(n5789), .Y(n4640) );
  CLKBUFX2 U4104 ( .A(n1052), .Y(n5789) );
  CLKINVX12 U4105 ( .A(n4671), .Y(n4641) );
  INVX8 U4106 ( .A(n4641), .Y(n4642) );
  INVX16 U4107 ( .A(n4641), .Y(n4643) );
  INVX4 U4108 ( .A(n5652), .Y(n6005) );
  NAND2X8 U4109 ( .A(cur_state), .B(n2662), .Y(n2661) );
  NOR2X2 U4110 ( .A(n6037), .B(n5660), .Y(n6034) );
  INVXL U4111 ( .A(n5652), .Y(n6037) );
  AOI221X4 U4112 ( .A0(n6623), .A1(n4696), .B0(n6558), .B1(n4649), .C0(n3769), 
        .Y(n3768) );
  INVX3 U4113 ( .A(n5788), .Y(n4644) );
  INVX8 U4114 ( .A(n4644), .Y(n4645) );
  CLKBUFX2 U4115 ( .A(n1052), .Y(n5788) );
  AOI221XL U4116 ( .A0(N3359), .A1(n3982), .B0(n5917), .B1(n3983), .C0(n4034), 
        .Y(n4029) );
  NOR2BX4 U4117 ( .AN(n5669), .B(n4696), .Y(n3983) );
  INVX3 U4118 ( .A(n5899), .Y(n4646) );
  CLKINVX12 U4119 ( .A(n4646), .Y(n4647) );
  INVXL U4120 ( .A(n5902), .Y(n5899) );
  CLKINVX8 U4121 ( .A(n5919), .Y(n5918) );
  INVX20 U4122 ( .A(n1050), .Y(n4648) );
  CLKINVX20 U4123 ( .A(n4648), .Y(n4649) );
  CLKINVX20 U4124 ( .A(n4648), .Y(n4650) );
  BUFX6 U4125 ( .A(n6291), .Y(n4651) );
  BUFX16 U4126 ( .A(n5774), .Y(n5773) );
  BUFX4 U4127 ( .A(n4804), .Y(n5774) );
  INVX3 U4128 ( .A(n5247), .Y(n4652) );
  INVX6 U4129 ( .A(n4652), .Y(n4653) );
  CLKINVX1 U4130 ( .A(n5663), .Y(n4654) );
  CLKINVX4 U4131 ( .A(n5663), .Y(n6226) );
  INVX1 U4132 ( .A(n5663), .Y(n6257) );
  CLKBUFX3 U4133 ( .A(n6257), .Y(n5740) );
  CLKBUFX6 U4134 ( .A(n5741), .Y(n5742) );
  MX4X4 U4135 ( .A(n5352), .B(n5342), .C(n5347), .D(n5337), .S0(N3334), .S1(
        N3333), .Y(N3364) );
  BUFX8 U4136 ( .A(N3364), .Y(n5663) );
  OAI22X2 U4137 ( .A0(n5913), .A1(n1810), .B0(n1823), .B1(n4637), .Y(n1822) );
  AOI221X2 U4138 ( .A0(N3358), .A1(n3982), .B0(n5921), .B1(n3983), .C0(n4026), 
        .Y(n4023) );
  NAND2X8 U4139 ( .A(cur_state), .B(n1567), .Y(n1566) );
  NAND2X8 U4140 ( .A(n5954), .B(n1788), .Y(n1787) );
  INVX4 U4141 ( .A(n1788), .Y(n6400) );
  AOI211X1 U4142 ( .A0(n6157), .A1(n6156), .B0(n6155), .C0(n6154), .Y(n6159)
         );
  NOR2BX1 U4143 ( .AN(n5653), .B(n5659), .Y(n6091) );
  AND2X4 U4144 ( .A(n4753), .B(n4032), .Y(n1058) );
  BUFX4 U4145 ( .A(n5970), .Y(n5057) );
  NOR2X1 U4146 ( .A(n6322), .B(n6333), .Y(n6334) );
  AND2X2 U4147 ( .A(n6233), .B(n6242), .Y(n6240) );
  INVX3 U4148 ( .A(n5931), .Y(n5930) );
  INVX2 U4149 ( .A(n5924), .Y(n5922) );
  INVX3 U4150 ( .A(n5939), .Y(n5936) );
  NOR2X1 U4151 ( .A(n6100), .B(n5652), .Y(n6096) );
  NOR2X1 U4152 ( .A(n6133), .B(n5660), .Y(n6129) );
  BUFX12 U4153 ( .A(n5962), .Y(n5961) );
  INVX1 U4154 ( .A(N3330), .Y(n5962) );
  AND3X4 U4155 ( .A(N5603), .B(N5602), .C(N5604), .Y(n4056) );
  OAI31X1 U4156 ( .A0(n6288), .A1(n6287), .A2(n6286), .B0(n6285), .Y(N5602) );
  CLKINVX6 U4157 ( .A(n4805), .Y(n4762) );
  NAND2X2 U4158 ( .A(n4799), .B(n6127), .Y(N5080) );
  NOR3BX2 U4159 ( .AN(N3334), .B(n6574), .C(n4800), .Y(n3413) );
  NOR3BX2 U4160 ( .AN(N3334), .B(n6574), .C(n5958), .Y(n3730) );
  MX4X1 U4161 ( .A(n5502), .B(n5500), .C(n5501), .D(n5499), .S0(n5648), .S1(
        n5647), .Y(n5503) );
  MX4X1 U4162 ( .A(n4938), .B(n4936), .C(n4937), .D(n4935), .S0(n5068), .S1(
        n5969), .Y(n4939) );
  MX4X1 U4163 ( .A(n4948), .B(n4946), .C(n4947), .D(n4945), .S0(n5068), .S1(
        n5969), .Y(n4949) );
  CLKBUFX8 U4164 ( .A(N3331), .Y(n5959) );
  AOI221X1 U4165 ( .A0(n6603), .A1(n4696), .B0(n6538), .B1(n4650), .C0(n2618), 
        .Y(n2617) );
  OAI22X1 U4166 ( .A0(n5913), .A1(n1932), .B0(n1944), .B1(n4637), .Y(n1943) );
  AOI221XL U4167 ( .A0(n6614), .A1(n4696), .B0(n6549), .B1(n4650), .C0(n1603), 
        .Y(n1602) );
  AOI221X1 U4168 ( .A0(n6597), .A1(n4696), .B0(n6532), .B1(n4649), .C0(n2024), 
        .Y(n2023) );
  NAND4X2 U4169 ( .A(n5667), .B(n6663), .C(n6664), .D(n6659), .Y(n1041) );
  MX4X1 U4170 ( .A(n5472), .B(n5470), .C(n5471), .D(n5469), .S0(n5649), .S1(
        n5647), .Y(n5473) );
  BUFX4 U4171 ( .A(n5457), .Y(N3375) );
  CLKBUFX8 U4172 ( .A(N3354), .Y(n5659) );
  OAI22X2 U4173 ( .A0(n5916), .A1(n3480), .B0(n3490), .B1(n4637), .Y(n3489) );
  OAI22X2 U4174 ( .A0(n5912), .A1(n3319), .B0(n3329), .B1(n4637), .Y(n3328) );
  INVX6 U4175 ( .A(n3852), .Y(n6349) );
  OAI22X2 U4176 ( .A0(n5913), .A1(n3358), .B0(n3368), .B1(n4637), .Y(n3367) );
  INVX6 U4177 ( .A(n4874), .Y(n2823) );
  OAI22X2 U4178 ( .A0(n5912), .A1(n3397), .B0(n3408), .B1(n4637), .Y(n3407) );
  OAI22X2 U4179 ( .A0(n5912), .A1(n3241), .B0(n3251), .B1(n4637), .Y(n3250) );
  OAI22X2 U4180 ( .A0(n5915), .A1(n2924), .B0(n2934), .B1(n4637), .Y(n2933) );
  OAI22X2 U4181 ( .A0(n5915), .A1(n3202), .B0(n3212), .B1(n4637), .Y(n3211) );
  INVX6 U4182 ( .A(n4873), .Y(n2862) );
  OAI22X2 U4183 ( .A0(n5912), .A1(n3441), .B0(n3451), .B1(n4637), .Y(n3450) );
  OAI22X2 U4184 ( .A0(n5913), .A1(n3280), .B0(n3290), .B1(n4637), .Y(n3289) );
  NAND2BX1 U4185 ( .AN(N3357), .B(n5926), .Y(n6302) );
  NOR2BX2 U4186 ( .AN(N3355), .B(n5936), .Y(n6150) );
  NOR2X1 U4187 ( .A(n6265), .B(n6277), .Y(n6278) );
  NOR2X1 U4188 ( .A(n6107), .B(n6119), .Y(n6120) );
  NOR3BX1 U4189 ( .AN(n6339), .B(n6338), .C(n6324), .Y(n6325) );
  NOR2X1 U4190 ( .A(n5979), .B(n5991), .Y(n5992) );
  INVX3 U4191 ( .A(N3323), .Y(n5967) );
  BUFX12 U4192 ( .A(n5967), .Y(n5965) );
  AOI211X1 U4193 ( .A0(n6202), .A1(n6214), .B0(n6201), .C0(n6217), .Y(n6203)
         );
  CLKINVX1 U4194 ( .A(n6237), .Y(n6259) );
  AOI211X1 U4195 ( .A0(n6171), .A1(n6183), .B0(n6170), .C0(n6186), .Y(n6172)
         );
  AOI31X1 U4196 ( .A0(n6026), .A1(n6011), .A2(n6010), .B0(n6023), .Y(n6013) );
  OAI211X1 U4197 ( .A0(n6009), .A1(n6036), .B0(n6008), .C0(n6018), .Y(n6010)
         );
  NOR2X1 U4198 ( .A(n6012), .B(n6024), .Y(n6025) );
  NAND2BX1 U4199 ( .AN(n6034), .B(n6016), .Y(n6029) );
  NAND2BX1 U4200 ( .AN(n6001), .B(n5983), .Y(n5996) );
  NAND3X1 U4201 ( .A(n4790), .B(n4791), .C(n4676), .Y(n4792) );
  NAND3X1 U4202 ( .A(n4767), .B(n4768), .C(n4769), .Y(n4770) );
  NAND3X1 U4203 ( .A(n4796), .B(n4797), .C(n4798), .Y(n4799) );
  CLKINVX1 U4204 ( .A(n6128), .Y(n4798) );
  INVX3 U4205 ( .A(n6078), .Y(n6102) );
  CLKINVX1 U4206 ( .A(N3321), .Y(n6499) );
  CLKINVX1 U4207 ( .A(N3320), .Y(n5968) );
  INVX6 U4208 ( .A(n4032), .Y(n6416) );
  CLKBUFX3 U4209 ( .A(n5445), .Y(n5446) );
  OAI22XL U4210 ( .A0(n3980), .A1(n5684), .B0(n3981), .B1(n5737), .Y(n4007) );
  NAND2BX2 U4211 ( .AN(N3324), .B(n5082), .Y(\sub_80/carry[2] ) );
  NOR2X1 U4212 ( .A(n5971), .B(n5963), .Y(n5972) );
  MX4X1 U4213 ( .A(n5567), .B(n5565), .C(n5566), .D(n5564), .S0(n5648), .S1(
        n5267), .Y(n5568) );
  NOR3BX2 U4214 ( .AN(n5963), .B(n5964), .C(n5634), .Y(n1739) );
  NOR3BX2 U4215 ( .AN(n5963), .B(n5964), .C(n5631), .Y(n1740) );
  NOR3BX2 U4216 ( .AN(n5969), .B(n4635), .C(n5634), .Y(n1782) );
  NOR3BX2 U4217 ( .AN(n5959), .B(n5961), .C(N3323), .Y(n1783) );
  NOR3BX2 U4218 ( .AN(N3334), .B(n5958), .C(N3333), .Y(n3096) );
  NOR3X2 U4219 ( .A(n5252), .B(n5963), .C(n5964), .Y(n1563) );
  NOR3X2 U4220 ( .A(n4749), .B(n5963), .C(n5634), .Y(n1064) );
  NOR3BX2 U4221 ( .AN(n5963), .B(n5634), .C(n4749), .Y(n1651) );
  NOR3BX2 U4222 ( .AN(n5963), .B(n5634), .C(n4749), .Y(n1652) );
  NOR3X2 U4223 ( .A(n5966), .B(n5963), .C(n5964), .Y(n1607) );
  NOR3X2 U4224 ( .A(n5252), .B(n5969), .C(n4634), .Y(n1605) );
  NOR3BX2 U4225 ( .AN(N3322), .B(n6499), .C(n5968), .Y(n3729) );
  NOR3BX2 U4226 ( .AN(n5673), .B(n6666), .C(n5955), .Y(n3415) );
  NOR3BX2 U4227 ( .AN(N3322), .B(n6499), .C(N3320), .Y(n3412) );
  NOR3BX2 U4228 ( .AN(n5673), .B(n4893), .C(N3339), .Y(n3098) );
  NOR3BX2 U4229 ( .AN(N3322), .B(n5968), .C(N3321), .Y(n3095) );
  NOR3BX2 U4230 ( .AN(N3334), .B(n4800), .C(N3333), .Y(n2779) );
  NOR3BX2 U4231 ( .AN(n5673), .B(n5955), .C(N3339), .Y(n2781) );
  NOR3BX2 U4232 ( .AN(N3322), .B(N3320), .C(N3321), .Y(n2778) );
  NOR3X2 U4233 ( .A(n5968), .B(N3322), .C(n6499), .Y(n2461) );
  NOR3X2 U4234 ( .A(N3320), .B(N3322), .C(n6499), .Y(n2144) );
  NOR3X2 U4235 ( .A(N3321), .B(N3322), .C(n5968), .Y(n1826) );
  NOR3X2 U4236 ( .A(n5674), .B(n5673), .C(n4893), .Y(n1829) );
  NOR3BX2 U4237 ( .AN(n5959), .B(n5634), .C(n5960), .Y(n1694) );
  NOR3BX2 U4238 ( .AN(n5969), .B(n5634), .C(n5058), .Y(n1693) );
  NOR3X2 U4239 ( .A(n4749), .B(n5963), .C(n5966), .Y(n1519) );
  NOR3X2 U4240 ( .A(n5063), .B(n5969), .C(n5634), .Y(n1517) );
  NOR3X2 U4241 ( .A(N3321), .B(N3322), .C(N3320), .Y(n1059) );
  NOR3X2 U4242 ( .A(n5674), .B(n5673), .C(n5955), .Y(n1065) );
  CLKBUFX16 U4243 ( .A(n1049), .Y(n4696) );
  INVX12 U4244 ( .A(n4825), .Y(n1050) );
  MX4X1 U4245 ( .A(n5216), .B(n5214), .C(n5215), .D(n5213), .S0(n5270), .S1(
        n5268), .Y(n5217) );
  OAI22XL U4246 ( .A0(n3980), .A1(n5699), .B0(n3981), .B1(n5750), .Y(n4031) );
  MX4X1 U4247 ( .A(\img_buff[28][2] ), .B(\img_buff[29][2] ), .C(
        \img_buff[30][2] ), .D(\img_buff[31][2] ), .S0(n5435), .S1(n4699), .Y(
        n5323) );
  MX4X1 U4248 ( .A(\img_buff[20][2] ), .B(\img_buff[21][2] ), .C(
        \img_buff[22][2] ), .D(\img_buff[23][2] ), .S0(n5435), .S1(n4699), .Y(
        n5325) );
  MX4X1 U4249 ( .A(\img_buff[12][2] ), .B(\img_buff[13][2] ), .C(
        \img_buff[14][2] ), .D(\img_buff[15][2] ), .S0(n5435), .S1(n4699), .Y(
        n5328) );
  MX4X1 U4250 ( .A(\img_buff[36][2] ), .B(\img_buff[37][2] ), .C(
        \img_buff[38][2] ), .D(\img_buff[39][2] ), .S0(n5435), .S1(n4699), .Y(
        n5320) );
  MX4X1 U4251 ( .A(\img_buff[44][2] ), .B(\img_buff[45][2] ), .C(
        \img_buff[46][2] ), .D(\img_buff[47][2] ), .S0(n5245), .S1(n5641), .Y(
        n5509) );
  AOI221X1 U4252 ( .A0(N3357), .A1(n3977), .B0(n5925), .B1(n3978), .C0(n4019), 
        .Y(n4018) );
  MX4X1 U4253 ( .A(n5562), .B(n5560), .C(n5561), .D(n5559), .S0(n5649), .S1(
        n5963), .Y(n5563) );
  MX4X1 U4254 ( .A(n5557), .B(n5555), .C(n5556), .D(n5554), .S0(n5648), .S1(
        n5269), .Y(n5558) );
  MX4X1 U4255 ( .A(n5527), .B(n5525), .C(n5526), .D(n5524), .S0(n5648), .S1(
        n5963), .Y(n5528) );
  OA22X1 U4256 ( .A0(n1032), .A1(n5772), .B0(n5771), .B1(n1033), .Y(n1056) );
  AOI221X1 U4257 ( .A0(n6584), .A1(n4696), .B0(n6519), .B1(n4650), .C0(n3647), 
        .Y(n3646) );
  OAI221XL U4258 ( .A0(n5780), .A1(n3635), .B0(n4665), .B1(n3648), .C0(n3649), 
        .Y(n3644) );
  OA22X1 U4259 ( .A0(n3486), .A1(n5773), .B0(n5767), .B1(n3480), .Y(n3493) );
  OA22X1 U4260 ( .A0(n3325), .A1(n5773), .B0(n5767), .B1(n3319), .Y(n3332) );
  AOI221X1 U4261 ( .A0(n6586), .A1(n4696), .B0(n6521), .B1(n4650), .C0(n3013), 
        .Y(n3012) );
  OA22X1 U4262 ( .A0(n3008), .A1(n5772), .B0(n5768), .B1(n3002), .Y(n3015) );
  OA22X1 U4263 ( .A0(n2535), .A1(n5773), .B0(n5769), .B1(n2529), .Y(n2542) );
  OA22X1 U4264 ( .A0(n2374), .A1(n5773), .B0(n5769), .B1(n2368), .Y(n2381) );
  OA22X1 U4265 ( .A0(n2218), .A1(n5773), .B0(n5769), .B1(n2212), .Y(n2225) );
  AOI221X1 U4266 ( .A0(n6589), .A1(n4696), .B0(n6524), .B1(n4650), .C0(n2062), 
        .Y(n2061) );
  OAI22XL U4267 ( .A0(n4640), .A1(n2051), .B0(n5785), .B1(n2057), .Y(n2062) );
  OAI221XL U4268 ( .A0(n5778), .A1(n2050), .B0(n4661), .B1(n2063), .C0(n2064), 
        .Y(n2059) );
  OA22X1 U4269 ( .A0(n2057), .A1(n5773), .B0(n5770), .B1(n2051), .Y(n2064) );
  NAND2X1 U4270 ( .A(n1737), .B(n1059), .Y(n1721) );
  AOI221X1 U4271 ( .A0(n6600), .A1(n4696), .B0(n6535), .B1(n4650), .C0(n3569), 
        .Y(n3568) );
  OAI221XL U4272 ( .A0(n5780), .A1(n3557), .B0(n4664), .B1(n3570), .C0(n3571), 
        .Y(n3566) );
  AND3X2 U4273 ( .A(n4775), .B(n4776), .C(n4670), .Y(n4051) );
  OA22X1 U4274 ( .A0(n4047), .A1(n5772), .B0(n5767), .B1(n4041), .Y(n4055) );
  OA22X1 U4275 ( .A0(n3525), .A1(n5773), .B0(n5767), .B1(n3519), .Y(n3532) );
  AOI221X1 U4276 ( .A0(n6608), .A1(n4696), .B0(n6543), .B1(n4650), .C0(n3530), 
        .Y(n3529) );
  OA22X1 U4277 ( .A0(n3364), .A1(n5773), .B0(n5767), .B1(n3358), .Y(n3371) );
  AOI221X1 U4278 ( .A0(n6578), .A1(n4696), .B0(n6513), .B1(n4650), .C0(n3052), 
        .Y(n3051) );
  OA22X1 U4279 ( .A0(n3047), .A1(n5772), .B0(n5768), .B1(n3041), .Y(n3054) );
  OAI221XL U4280 ( .A0(n5779), .A1(n2723), .B0(n4657), .B1(n2736), .C0(n2737), 
        .Y(n2732) );
  OA22X1 U4281 ( .A0(n2730), .A1(n5773), .B0(n5768), .B1(n2724), .Y(n2737) );
  OA22X1 U4282 ( .A0(n2574), .A1(n5773), .B0(n5769), .B1(n2568), .Y(n2581) );
  OA22X1 U4283 ( .A0(n2413), .A1(n5773), .B0(n5769), .B1(n2407), .Y(n2420) );
  AOI221X1 U4284 ( .A0(n6581), .A1(n4696), .B0(n6516), .B1(n4650), .C0(n2101), 
        .Y(n2100) );
  OAI22XL U4285 ( .A0(n4640), .A1(n2090), .B0(n5785), .B1(n2096), .Y(n2101) );
  OA22X1 U4286 ( .A0(n2096), .A1(n5773), .B0(n5770), .B1(n2090), .Y(n2103) );
  NAND2X1 U4287 ( .A(n1782), .B(n1059), .Y(n1765) );
  OA22X1 U4288 ( .A0(n1769), .A1(n5772), .B0(n5770), .B1(n1765), .Y(n1781) );
  AOI221X1 U4289 ( .A0(n6592), .A1(n4696), .B0(n6527), .B1(n4650), .C0(n3608), 
        .Y(n3607) );
  OAI221XL U4290 ( .A0(n5780), .A1(n3596), .B0(n4665), .B1(n3609), .C0(n3610), 
        .Y(n3605) );
  BUFX8 U4291 ( .A(N3361), .Y(n5660) );
  BUFX4 U4292 ( .A(N3345), .Y(n5652) );
  MX4X1 U4293 ( .A(n5034), .B(n5024), .C(n5029), .D(n5019), .S0(N3322), .S1(
        N3321), .Y(N3345) );
  OA22X1 U4294 ( .A0(n2652), .A1(n5773), .B0(n5768), .B1(n2646), .Y(n2659) );
  OA22X1 U4295 ( .A0(n2335), .A1(n5773), .B0(n5769), .B1(n2329), .Y(n2342) );
  INVX3 U4296 ( .A(N3369), .Y(n5947) );
  CLKBUFX3 U4297 ( .A(n5463), .Y(N3369) );
  AOI221X1 U4298 ( .A0(n6617), .A1(n4696), .B0(n6552), .B1(n4650), .C0(n3174), 
        .Y(n3173) );
  OA22X1 U4299 ( .A0(n1897), .A1(n5772), .B0(n5770), .B1(n1893), .Y(n1907) );
  AOI221X1 U4300 ( .A0(n6621), .A1(n4696), .B0(n6556), .B1(n4650), .C0(n1906), 
        .Y(n1905) );
  NAND2X1 U4301 ( .A(n1826), .B(n1561), .Y(n1893) );
  OA22X1 U4302 ( .A0(n3403), .A1(n5773), .B0(n5767), .B1(n3397), .Y(n3411) );
  OAI221XL U4303 ( .A0(n5779), .A1(n3240), .B0(n4659), .B1(n3253), .C0(n3254), 
        .Y(n3249) );
  OAI221XL U4304 ( .A0(n5779), .A1(n3079), .B0(n4660), .B1(n3093), .C0(n3094), 
        .Y(n3089) );
  OA22X1 U4305 ( .A0(n2930), .A1(n5773), .B0(n5768), .B1(n2924), .Y(n2937) );
  OA22X1 U4306 ( .A0(n2769), .A1(n5773), .B0(n5768), .B1(n2763), .Y(n2777) );
  AOI221X1 U4307 ( .A0(n6636), .A1(n4696), .B0(n6571), .B1(n4650), .C0(n2141), 
        .Y(n2140) );
  OAI22XL U4308 ( .A0(n4640), .A1(n2129), .B0(n5785), .B1(n2135), .Y(n2141) );
  OA22X1 U4309 ( .A0(n2135), .A1(n5772), .B0(n5769), .B1(n2129), .Y(n2143) );
  AOI221X1 U4310 ( .A0(n6605), .A1(n4696), .B0(n6540), .B1(n4650), .C0(n1984), 
        .Y(n1983) );
  OAI22XL U4311 ( .A0(n4639), .A1(n1971), .B0(n5785), .B1(n1975), .Y(n1984) );
  OA22X1 U4312 ( .A0(n1975), .A1(n5772), .B0(n5770), .B1(n1971), .Y(n1985) );
  NAND2X1 U4313 ( .A(n1826), .B(n1060), .Y(n1810) );
  NAND2X1 U4314 ( .A(n1649), .B(n1059), .Y(n1633) );
  OA22X1 U4315 ( .A0(n3208), .A1(n5773), .B0(n5767), .B1(n3202), .Y(n3215) );
  NAND2X1 U4316 ( .A(n1826), .B(n1605), .Y(n1932) );
  OA22X1 U4317 ( .A0(n3447), .A1(n5773), .B0(n5767), .B1(n3441), .Y(n3454) );
  OA22X1 U4318 ( .A0(n3286), .A1(n5773), .B0(n5767), .B1(n3280), .Y(n3293) );
  OAI221XL U4319 ( .A0(n5779), .A1(n3123), .B0(n4658), .B1(n3136), .C0(n3137), 
        .Y(n3132) );
  OA22X1 U4320 ( .A0(n2969), .A1(n5772), .B0(n5768), .B1(n2963), .Y(n2976) );
  OAI22X1 U4321 ( .A0(n4645), .A1(n2963), .B0(n5785), .B1(n2969), .Y(n2974) );
  OA22X1 U4322 ( .A0(n2813), .A1(n5773), .B0(n5768), .B1(n2807), .Y(n2820) );
  OA22X1 U4323 ( .A0(n2496), .A1(n5773), .B0(n5769), .B1(n2490), .Y(n2503) );
  OA22X1 U4324 ( .A0(n2179), .A1(n5773), .B0(n5769), .B1(n2173), .Y(n2186) );
  NAND2X1 U4325 ( .A(n1826), .B(n1517), .Y(n1854) );
  OA22X1 U4326 ( .A0(n1858), .A1(n4804), .B0(n5770), .B1(n1854), .Y(n1868) );
  NAND2X1 U4327 ( .A(n1693), .B(n1059), .Y(n1677) );
  AOI211X1 U4328 ( .A0(n5934), .A1(n6483), .B0(n1797), .C0(n5889), .Y(n1796)
         );
  INVX6 U4329 ( .A(n4824), .Y(N3359) );
  INVX6 U4330 ( .A(n4815), .Y(N3351) );
  MX4X2 U4331 ( .A(n4934), .B(n4924), .C(n4929), .D(n4919), .S0(N3322), .S1(
        N3321), .Y(N3350) );
  MX4X1 U4332 ( .A(n5492), .B(n5490), .C(n5491), .D(n5489), .S0(n5649), .S1(
        n5267), .Y(n5493) );
  MX4X1 U4333 ( .A(n5487), .B(n5485), .C(n5486), .D(n5484), .S0(n5649), .S1(
        n5267), .Y(n5488) );
  BUFX12 U4334 ( .A(N3349), .Y(n5656) );
  MX4X1 U4335 ( .A(n4953), .B(n4951), .C(n4952), .D(n4950), .S0(n5068), .S1(
        n5969), .Y(n4954) );
  INVX6 U4336 ( .A(n4808), .Y(N3357) );
  INVX4 U4337 ( .A(n5459), .Y(n5927) );
  BUFX8 U4338 ( .A(N3363), .Y(n5662) );
  MX4X2 U4339 ( .A(n5372), .B(n5362), .C(n5367), .D(n5357), .S0(N3334), .S1(
        N3333), .Y(N3363) );
  MX4X1 U4340 ( .A(n5371), .B(n5369), .C(n5370), .D(n5368), .S0(n4800), .S1(
        n5456), .Y(n5372) );
  CLKINVX12 U4341 ( .A(n5927), .Y(n5926) );
  BUFX12 U4342 ( .A(N3362), .Y(n5661) );
  MX4X2 U4343 ( .A(n5392), .B(n5382), .C(n5387), .D(n5377), .S0(N3334), .S1(
        N3333), .Y(N3362) );
  BUFX4 U4344 ( .A(N3346), .Y(n5653) );
  MX4X1 U4345 ( .A(n5014), .B(n5004), .C(n5009), .D(n4999), .S0(N3322), .S1(
        N3321), .Y(N3346) );
  INVX3 U4346 ( .A(n997), .Y(n5902) );
  INVX3 U4347 ( .A(n4838), .Y(n2662) );
  AOI221X1 U4348 ( .A0(n2682), .A1(n4701), .B0(n4697), .B1(n2693), .C0(n2694), 
        .Y(n2692) );
  OAI22X2 U4349 ( .A0(n5915), .A1(n2685), .B0(n2695), .B1(n4637), .Y(n2694) );
  INVX4 U4350 ( .A(n4811), .Y(n1699) );
  OAI221XL U4351 ( .A0(n5777), .A1(n1720), .B0(n4659), .B1(n1727), .C0(n1736), 
        .Y(n1732) );
  INVX4 U4352 ( .A(n4840), .Y(n2584) );
  AOI221X1 U4353 ( .A0(n2604), .A1(n4701), .B0(n4697), .B1(n2615), .C0(n2616), 
        .Y(n2614) );
  OAI22X2 U4354 ( .A0(n5914), .A1(n2607), .B0(n2617), .B1(n4637), .Y(n2616) );
  INVX3 U4355 ( .A(n4848), .Y(n2267) );
  INVX3 U4356 ( .A(n4849), .Y(n2228) );
  INVX12 U4357 ( .A(n5931), .Y(n5929) );
  INVX3 U4358 ( .A(n4844), .Y(n2423) );
  INVX4 U4359 ( .A(n4833), .Y(n1788) );
  OA22X2 U4360 ( .A0(n1819), .A1(n4627), .B0(n1042), .B1(n1820), .Y(n4833) );
  INVX4 U4361 ( .A(n4812), .Y(n1611) );
  OAI221XL U4362 ( .A0(n5777), .A1(n1632), .B0(n4659), .B1(n1639), .C0(n1648), 
        .Y(n1644) );
  INVX4 U4363 ( .A(n4831), .Y(n1910) );
  INVX8 U4364 ( .A(n4834), .Y(n1567) );
  OAI221XL U4365 ( .A0(n5777), .A1(n1588), .B0(n4660), .B1(n1595), .C0(n1604), 
        .Y(n1600) );
  INVX6 U4366 ( .A(n4877), .Y(n3735) );
  OA22X2 U4367 ( .A0(n3765), .A1(n4627), .B0(n1511), .B1(n3722), .Y(n4877) );
  INVX4 U4368 ( .A(n4813), .Y(n1988) );
  OAI22X1 U4369 ( .A0(n5913), .A1(n2010), .B0(n2023), .B1(n4637), .Y(n2022) );
  INVX4 U4370 ( .A(n4810), .Y(n1655) );
  NAND3X1 U4371 ( .A(n4750), .B(n4751), .C(n4752), .Y(n4175) );
  NAND3X1 U4372 ( .A(n4764), .B(n4765), .C(n4766), .Y(n4155) );
  NAND3X1 U4373 ( .A(n4780), .B(n4781), .C(n4782), .Y(n4183) );
  OR2X1 U4374 ( .A(n1887), .B(n1870), .Y(n4781) );
  NAND3X1 U4375 ( .A(n4759), .B(n4760), .C(n4761), .Y(n4543) );
  OR2X1 U4376 ( .A(n6354), .B(n5857), .Y(n4759) );
  OR2X1 U4377 ( .A(n3669), .B(n3651), .Y(n4760) );
  NAND3X1 U4378 ( .A(n4777), .B(n4778), .C(n4779), .Y(n4174) );
  OR2X1 U4379 ( .A(n1846), .B(n1831), .Y(n4778) );
  OAI222XL U4380 ( .A0(n6347), .A1(n5855), .B0(n3947), .B1(n3929), .C0(n701), 
        .C1(n3930), .Y(n4599) );
  OAI222XL U4381 ( .A0(n6351), .A1(n5856), .B0(n3791), .B1(n3773), .C0(n669), 
        .C1(n3774), .Y(n4567) );
  OAI222XL U4382 ( .A0(n6355), .A1(n5855), .B0(n3630), .B1(n3612), .C0(n637), 
        .C1(n3613), .Y(n4535) );
  OAI222XL U4383 ( .A0(n6359), .A1(n5855), .B0(n3474), .B1(n3456), .C0(n605), 
        .C1(n3457), .Y(n4503) );
  OAI222XL U4384 ( .A0(n6363), .A1(n5855), .B0(n3313), .B1(n3295), .C0(n573), 
        .C1(n3296), .Y(n4471) );
  OAI222XL U4385 ( .A0(n6367), .A1(n5855), .B0(n3157), .B1(n3139), .C0(n541), 
        .C1(n4674), .Y(n4439) );
  OAI222XL U4386 ( .A0(n6371), .A1(n5856), .B0(n2996), .B1(n2978), .C0(n509), 
        .C1(n2979), .Y(n4407) );
  OAI222XL U4387 ( .A0(n6375), .A1(n5856), .B0(n2840), .B1(n2822), .C0(n477), 
        .C1(n2823), .Y(n4375) );
  OAI222XL U4388 ( .A0(n6367), .A1(n5893), .B0(n3149), .B1(n3139), .C0(n537), 
        .C1(n4674), .Y(n4435) );
  OAI222XL U4389 ( .A0(n6349), .A1(n5856), .B0(n3869), .B1(n3851), .C0(n685), 
        .C1(n3852), .Y(n4583) );
  OAI222XL U4390 ( .A0(n6353), .A1(n5856), .B0(n3708), .B1(n3690), .C0(n653), 
        .C1(n5670), .Y(n4551) );
  OAI222XL U4391 ( .A0(n6357), .A1(n5855), .B0(n3552), .B1(n3534), .C0(n621), 
        .C1(n3535), .Y(n4519) );
  OAI222XL U4392 ( .A0(n6361), .A1(n5855), .B0(n3391), .B1(n3373), .C0(n589), 
        .C1(n3374), .Y(n4487) );
  OAI222XL U4393 ( .A0(n6365), .A1(n5855), .B0(n3235), .B1(n3217), .C0(n557), 
        .C1(n3218), .Y(n4455) );
  OAI222XL U4394 ( .A0(n6369), .A1(n5855), .B0(n3074), .B1(n3056), .C0(n525), 
        .C1(n3057), .Y(n4423) );
  OAI222XL U4395 ( .A0(n6373), .A1(n5856), .B0(n2918), .B1(n2900), .C0(n493), 
        .C1(n2901), .Y(n4391) );
  OAI222XL U4396 ( .A0(n6350), .A1(n5855), .B0(n3830), .B1(n3812), .C0(n677), 
        .C1(n3813), .Y(n4575) );
  OAI222XL U4397 ( .A0(n6358), .A1(n5855), .B0(n3513), .B1(n3495), .C0(n613), 
        .C1(n3496), .Y(n4511) );
  OAI222XL U4398 ( .A0(n6362), .A1(n5855), .B0(n3352), .B1(n3334), .C0(n581), 
        .C1(n3335), .Y(n4479) );
  OAI222XL U4399 ( .A0(n6366), .A1(n5855), .B0(n3196), .B1(n3178), .C0(n549), 
        .C1(n3179), .Y(n4447) );
  OAI222XL U4400 ( .A0(n6370), .A1(n5856), .B0(n3035), .B1(n3017), .C0(n517), 
        .C1(n3018), .Y(n4415) );
  OAI222XL U4401 ( .A0(n6374), .A1(n5856), .B0(n2879), .B1(n2861), .C0(n485), 
        .C1(n2862), .Y(n4383) );
  OAI222XL U4402 ( .A0(n6382), .A1(n5857), .B0(n2562), .B1(n2544), .C0(n421), 
        .C1(n2545), .Y(n4319) );
  OAI222XL U4403 ( .A0(n6401), .A1(n5858), .B0(n1759), .B1(n1742), .C0(n261), 
        .C1(n1743), .Y(n4159) );
  OAI222XL U4404 ( .A0(n3968), .A1(n5895), .B0(n4003), .B1(n3970), .C0(n705), 
        .C1(n6346), .Y(n4603) );
  OAI222XL U4405 ( .A0(n6348), .A1(n5857), .B0(n3908), .B1(n3890), .C0(n693), 
        .C1(n3891), .Y(n4591) );
  OAI222XL U4406 ( .A0(n6356), .A1(n5856), .B0(n3591), .B1(n3573), .C0(n629), 
        .C1(n3574), .Y(n4527) );
  OAI222XL U4407 ( .A0(n6360), .A1(n5855), .B0(n3435), .B1(n3417), .C0(n597), 
        .C1(n3418), .Y(n4495) );
  OAI222XL U4408 ( .A0(n6364), .A1(n5855), .B0(n3274), .B1(n3256), .C0(n565), 
        .C1(n3257), .Y(n4463) );
  OAI222XL U4409 ( .A0(n6368), .A1(n5855), .B0(n3118), .B1(n3100), .C0(n533), 
        .C1(n3101), .Y(n4431) );
  OAI222XL U4410 ( .A0(n6372), .A1(n5856), .B0(n2957), .B1(n2939), .C0(n501), 
        .C1(n4675), .Y(n4399) );
  OAI222XL U4411 ( .A0(n6372), .A1(n5894), .B0(n2949), .B1(n2939), .C0(n497), 
        .C1(n4675), .Y(n4395) );
  OAI222XL U4412 ( .A0(n6399), .A1(n5875), .B0(n1844), .B1(n1831), .C0(n275), 
        .C1(n4643), .Y(n4173) );
  NAND3XL U4413 ( .A(cmd_reg[2]), .B(n4060), .C(cmd_reg[1]), .Y(n972) );
  NAND2X8 U4414 ( .A(n5954), .B(n3735), .Y(n3734) );
  BUFX4 U4415 ( .A(n5245), .Y(n5251) );
  BUFX2 U4416 ( .A(n5254), .Y(n5244) );
  INVX4 U4417 ( .A(n5795), .Y(n5792) );
  CLKBUFX3 U4418 ( .A(n5775), .Y(n4655) );
  CLKBUFX3 U4419 ( .A(n4826), .Y(n4656) );
  INVX3 U4420 ( .A(n4656), .Y(n4657) );
  INVX3 U4421 ( .A(n4656), .Y(n4658) );
  INVX3 U4422 ( .A(n4656), .Y(n4659) );
  INVX3 U4423 ( .A(n4656), .Y(n4660) );
  INVX3 U4424 ( .A(n4656), .Y(n4661) );
  INVX3 U4425 ( .A(n4655), .Y(n4662) );
  INVX3 U4426 ( .A(n4662), .Y(n4663) );
  INVX3 U4427 ( .A(n4662), .Y(n4664) );
  INVX3 U4428 ( .A(n4662), .Y(n4665) );
  CLKINVX1 U4429 ( .A(n4826), .Y(n1055) );
  AO21X2 U4430 ( .A0(n4056), .A1(n5777), .B0(n6416), .Y(n4826) );
  INVX4 U4431 ( .A(n5763), .Y(n5758) );
  INVX4 U4432 ( .A(n5761), .Y(n5760) );
  INVX4 U4433 ( .A(n5762), .Y(n5759) );
  AOI211XL U4434 ( .A0(n5457), .A1(n6491), .B0(n1628), .C0(n5794), .Y(n1627)
         );
  AOI211XL U4435 ( .A0(n5457), .A1(n2546), .B0(n2563), .C0(n5792), .Y(n2562)
         );
  INVX3 U4436 ( .A(n5958), .Y(n5957) );
  CLKINVX6 U4437 ( .A(n5958), .Y(n4800) );
  OAI21X1 U4438 ( .A0(n4056), .A1(n4033), .B0(n4032), .Y(n4804) );
  OAI21X1 U4439 ( .A0(n4056), .A1(n4033), .B0(n4032), .Y(n4753) );
  CLKBUFX4 U4440 ( .A(n4753), .Y(n5772) );
  MX4X4 U4441 ( .A(n5523), .B(n5513), .C(n5518), .D(n5508), .S0(n5672), .S1(
        n5674), .Y(n5459) );
  MX4X1 U4442 ( .A(n4993), .B(n4991), .C(n4992), .D(n4990), .S0(n5067), .S1(
        n5066), .Y(n4994) );
  CLKBUFX3 U4443 ( .A(n5969), .Y(n5066) );
  NOR2BX2 U4444 ( .AN(N3351), .B(N3375), .Y(n6262) );
  INVX8 U4445 ( .A(n1007), .Y(n5882) );
  AOI221X1 U4446 ( .A0(N3355), .A1(n3977), .B0(n5935), .B1(n3978), .C0(n4007), 
        .Y(n4006) );
  AOI221X4 U4447 ( .A0(N3358), .A1(n3977), .B0(n5921), .B1(n3978), .C0(n4025), 
        .Y(n4024) );
  AOI221XL U4448 ( .A0(n5658), .A1(n3977), .B0(n5948), .B1(n3978), .C0(n3979), 
        .Y(n3976) );
  AOI221X1 U4449 ( .A0(N3359), .A1(n3977), .B0(n5917), .B1(n3978), .C0(n4031), 
        .Y(n4030) );
  AOI221X1 U4450 ( .A0(N3353), .A1(n3977), .B0(n5944), .B1(n3978), .C0(n3994), 
        .Y(n3993) );
  AOI221XL U4451 ( .A0(n4667), .A1(n3977), .B0(n5929), .B1(n3978), .C0(n4013), 
        .Y(n4012) );
  AOI221X1 U4452 ( .A0(n5659), .A1(n3977), .B0(n5941), .B1(n3978), .C0(n4001), 
        .Y(n3999) );
  CLKBUFX3 U4453 ( .A(N3324), .Y(n5266) );
  CLKINVX3 U4454 ( .A(n5824), .Y(n5816) );
  CLKINVX3 U4455 ( .A(n5826), .Y(n5817) );
  BUFX12 U4456 ( .A(n5076), .Y(n5436) );
  CLKBUFX6 U4457 ( .A(n5442), .Y(n5435) );
  CLKBUFX6 U4458 ( .A(n5626), .Y(n5629) );
  BUFX4 U4459 ( .A(n5970), .Y(n5056) );
  CLKBUFX3 U4460 ( .A(N3324), .Y(n5638) );
  XNOR2X4 U4461 ( .A(n4822), .B(n4823), .Y(n4666) );
  INVX16 U4462 ( .A(n4763), .Y(n5970) );
  MX4X4 U4463 ( .A(n5162), .B(n5152), .C(n5157), .D(n5147), .S0(n4666), .S1(
        N3327), .Y(n4667) );
  INVX6 U4464 ( .A(n4817), .Y(N3358) );
  MX4X2 U4465 ( .A(n5222), .B(n5212), .C(n5217), .D(n5207), .S0(n4666), .S1(
        N3327), .Y(N3353) );
  BUFX4 U4466 ( .A(n5650), .Y(n5648) );
  CLKINVX1 U4467 ( .A(n5655), .Y(n6067) );
  BUFX4 U4468 ( .A(n5057), .Y(n5059) );
  MXI4X2 U4469 ( .A(n5102), .B(n5092), .C(n5097), .D(n5087), .S0(n4666), .S1(
        N3327), .Y(n4824) );
  BUFX12 U4470 ( .A(n5449), .Y(n4699) );
  INVX1 U4471 ( .A(n5655), .Y(n6004) );
  CLKINVX1 U4472 ( .A(n5666), .Y(n6509) );
  CLKBUFX3 U4473 ( .A(n6507), .Y(n5743) );
  CLKBUFX3 U4474 ( .A(n5963), .Y(n5269) );
  INVX1 U4475 ( .A(n5652), .Y(n6068) );
  CLKBUFX2 U4476 ( .A(n5445), .Y(n5449) );
  BUFX4 U4477 ( .A(n5064), .Y(n5061) );
  BUFX4 U4478 ( .A(n5057), .Y(n5058) );
  MXI4X2 U4479 ( .A(n5122), .B(n5112), .C(n5117), .D(n5107), .S0(n4666), .S1(
        N3327), .Y(n4817) );
  INVX3 U4480 ( .A(N3338), .Y(n5956) );
  INVX1 U4481 ( .A(n5665), .Y(n6225) );
  CLKBUFX6 U4482 ( .A(N3344), .Y(n5651) );
  CLKINVX12 U4483 ( .A(n5961), .Y(n5960) );
  INVX1 U4484 ( .A(n5653), .Y(n6418) );
  BUFX4 U4485 ( .A(n5056), .Y(n5062) );
  CLKBUFX6 U4486 ( .A(n5637), .Y(n5626) );
  CLKINVX3 U4487 ( .A(n5862), .Y(n5860) );
  CLKINVX3 U4488 ( .A(n5862), .Y(n5861) );
  CLKBUFX3 U4489 ( .A(N3324), .Y(n5256) );
  INVX1 U4490 ( .A(n5652), .Y(n6417) );
  INVX1 U4491 ( .A(n5657), .Y(n6422) );
  INVX1 U4492 ( .A(n5655), .Y(n6420) );
  INVX1 U4493 ( .A(n5662), .Y(n6506) );
  CLKBUFX3 U4494 ( .A(n5731), .Y(n5730) );
  INVX1 U4495 ( .A(n5660), .Y(n6504) );
  INVXL U4496 ( .A(n5656), .Y(n6421) );
  INVXL U4497 ( .A(n5654), .Y(n6419) );
  CLKBUFX2 U4498 ( .A(n4815), .Y(n5698) );
  CLKBUFX2 U4499 ( .A(n4816), .Y(n5711) );
  BUFX4 U4500 ( .A(N3320), .Y(n5068) );
  CLKBUFX6 U4501 ( .A(N3319), .Y(n5969) );
  BUFX16 U4502 ( .A(N3325), .Y(n5963) );
  MXI4X1 U4503 ( .A(n5623), .B(n5613), .C(n5618), .D(n5608), .S0(n5672), .S1(
        n5674), .Y(n4668) );
  BUFX2 U4504 ( .A(N3323), .Y(n5255) );
  CLKBUFX3 U4505 ( .A(n6418), .Y(n5681) );
  INVX1 U4506 ( .A(n5665), .Y(n6508) );
  CLKBUFX2 U4507 ( .A(n976), .Y(n5912) );
  INVX6 U4508 ( .A(n4816), .Y(N3355) );
  MXI4X2 U4509 ( .A(n5182), .B(n5172), .C(n5177), .D(n5167), .S0(n4666), .S1(
        N3327), .Y(n4816) );
  INVX3 U4510 ( .A(n1002), .Y(n5892) );
  CLKXOR2X4 U4511 ( .A(n5955), .B(\sub_80/carry[3] ), .Y(N3320) );
  INVX1 U4512 ( .A(n5673), .Y(n4819) );
  OA22X2 U4513 ( .A0(n3974), .A1(n3975), .B0(n3976), .B1(n5668), .Y(n4669) );
  INVX3 U4514 ( .A(n5458), .Y(n5924) );
  OA22XL U4515 ( .A0(n5786), .A1(n4041), .B0(n5785), .B1(n4047), .Y(n4670) );
  CLKBUFX2 U4516 ( .A(n1054), .Y(n5776) );
  INVX3 U4517 ( .A(n5461), .Y(n5939) );
  CLKINVX1 U4518 ( .A(n5460), .Y(n5933) );
  CLKBUFX2 U4519 ( .A(n5963), .Y(n5647) );
  INVX3 U4520 ( .A(n1017), .Y(n5862) );
  BUFX16 U4521 ( .A(n5960), .Y(n5450) );
  CLKBUFX2 U4522 ( .A(n4668), .Y(n5950) );
  CLKBUFX2 U4523 ( .A(n5947), .Y(n5946) );
  INVX6 U4524 ( .A(n5890), .Y(n5889) );
  INVX3 U4525 ( .A(n1012), .Y(n5871) );
  INVX3 U4526 ( .A(n5862), .Y(n5859) );
  OAI22X4 U4527 ( .A0(n1863), .A1(n4627), .B0(n1511), .B1(n1820), .Y(n4671) );
  OA22X2 U4528 ( .A0(n3992), .A1(n3975), .B0(n3993), .B1(n5668), .Y(n4814) );
  OR3X2 U4529 ( .A(n4801), .B(n4802), .C(n4803), .Y(n4672) );
  OA21X2 U4530 ( .A0(n5972), .A1(n5956), .B0(n5973), .Y(n4673) );
  OAI22X4 U4531 ( .A0(n3170), .A1(n4627), .B0(n1555), .B1(n3088), .Y(n4674) );
  OAI22X4 U4532 ( .A0(n2970), .A1(n4627), .B0(n1687), .B1(n2771), .Y(n4675) );
  BUFX4 U4533 ( .A(n5960), .Y(n5455) );
  BUFX4 U4534 ( .A(n5455), .Y(n5445) );
  CLKBUFX3 U4535 ( .A(n5445), .Y(n5447) );
  OR2X1 U4536 ( .A(n4786), .B(n6091), .Y(n4676) );
  MX4X1 U4537 ( .A(n5563), .B(n5553), .C(n5558), .D(n5548), .S0(n5672), .S1(
        n5674), .Y(n5461) );
  MX4X1 U4538 ( .A(n5503), .B(n5493), .C(n5498), .D(n5488), .S0(n5672), .S1(
        n5674), .Y(n5458) );
  CLKBUFX3 U4539 ( .A(n5776), .Y(n5780) );
  INVX12 U4540 ( .A(n5949), .Y(n5948) );
  INVX3 U4541 ( .A(n5462), .Y(n5943) );
  INVX4 U4542 ( .A(n5947), .Y(n5945) );
  INVX8 U4543 ( .A(n5947), .Y(n5944) );
  CLKBUFX6 U4544 ( .A(n5624), .Y(n5634) );
  AND2X1 U4545 ( .A(n1451), .B(n1436), .Y(n4677) );
  AND2X2 U4546 ( .A(n1451), .B(n1432), .Y(n4678) );
  AND2X2 U4547 ( .A(n1446), .B(n1434), .Y(n4679) );
  AND2X2 U4548 ( .A(n1446), .B(n1432), .Y(n4680) );
  AND2XL U4549 ( .A(n1446), .B(n1436), .Y(n4681) );
  AND2X2 U4550 ( .A(n1431), .B(n1441), .Y(n4682) );
  AND2X2 U4551 ( .A(n1432), .B(n1460), .Y(n4683) );
  AND2X2 U4552 ( .A(n1436), .B(n1460), .Y(n4684) );
  CLKINVX2 U4553 ( .A(n6691), .Y(n6655) );
  INVX3 U4554 ( .A(n4677), .Y(n4685) );
  NAND2X2 U4555 ( .A(n1436), .B(n1441), .Y(n1092) );
  INVX3 U4556 ( .A(n4681), .Y(n4686) );
  INVX3 U4557 ( .A(n4678), .Y(n4687) );
  INVX3 U4558 ( .A(n4680), .Y(n4688) );
  INVX3 U4559 ( .A(n4679), .Y(n4689) );
  INVX3 U4560 ( .A(n4684), .Y(n4690) );
  INVX3 U4561 ( .A(n4683), .Y(n4691) );
  INVX3 U4562 ( .A(n4682), .Y(n4692) );
  NOR3X2 U4563 ( .A(n5060), .B(n5969), .C(n5966), .Y(n1060) );
  NOR3X2 U4564 ( .A(n5966), .B(n5969), .C(n4633), .Y(n1561) );
  CLKBUFX3 U4565 ( .A(n5967), .Y(n5966) );
  INVXL U4566 ( .A(n4729), .Y(n4693) );
  INVX12 U4567 ( .A(n4693), .Y(busy) );
  CLKBUFX3 U4568 ( .A(n5966), .Y(n5437) );
  NAND2X4 U4569 ( .A(n5952), .B(n1479), .Y(n1478) );
  NAND2X4 U4570 ( .A(n5953), .B(n1523), .Y(n1522) );
  NOR2X1 U4571 ( .A(n5946), .B(n5660), .Y(n6343) );
  CLKBUFX2 U4572 ( .A(n5255), .Y(n5246) );
  AND2X2 U4573 ( .A(n6264), .B(n6274), .Y(n6271) );
  AOI221X1 U4574 ( .A0(n1630), .A1(n4701), .B0(n4697), .B1(n1644), .C0(n1645), 
        .Y(n1642) );
  AOI221X1 U4575 ( .A0(n1674), .A1(n4701), .B0(n4697), .B1(n1688), .C0(n1689), 
        .Y(n1686) );
  OAI221X1 U4576 ( .A0(n5777), .A1(n1676), .B0(n4664), .B1(n1683), .C0(n1692), 
        .Y(n1688) );
  AOI221X1 U4577 ( .A0(n1718), .A1(n4701), .B0(n4697), .B1(n1732), .C0(n1733), 
        .Y(n1730) );
  OAI31X4 U4578 ( .A0(n6256), .A1(n6255), .A2(n6254), .B0(n6253), .Y(N5343) );
  NOR2BX1 U4579 ( .AN(n5659), .B(n5941), .Y(n6309) );
  OAI31X1 U4580 ( .A0(n6344), .A1(n6343), .A2(n6342), .B0(n6341), .Y(N5604) );
  NAND2BX1 U4581 ( .AN(n6343), .B(n6326), .Y(n6338) );
  CLKINVX1 U4582 ( .A(N3375), .Y(n5919) );
  BUFX4 U4583 ( .A(n5056), .Y(n4695) );
  BUFX6 U4584 ( .A(n5970), .Y(n5064) );
  BUFX4 U4585 ( .A(n5064), .Y(n5060) );
  NAND2X2 U4586 ( .A(n4036), .B(n4035), .Y(n1049) );
  BUFX4 U4587 ( .A(n5256), .Y(n5641) );
  BUFX4 U4588 ( .A(n5441), .Y(n5076) );
  NOR3BX1 U4589 ( .AN(n6156), .B(n6155), .C(n6141), .Y(n6142) );
  AOI211X2 U4590 ( .A0(n6140), .A1(n6151), .B0(n6139), .C0(n6154), .Y(n6141)
         );
  CLKINVX12 U4591 ( .A(n3968), .Y(n6346) );
  MX4XL U4592 ( .A(\img_buff[4][2] ), .B(\img_buff[5][2] ), .C(
        \img_buff[6][2] ), .D(\img_buff[7][2] ), .S0(n5435), .S1(n5960), .Y(
        n5330) );
  INVX6 U4593 ( .A(n4643), .Y(n6399) );
  NAND2X8 U4594 ( .A(n5954), .B(n4642), .Y(n1831) );
  MX4X2 U4595 ( .A(n4963), .B(n4961), .C(n4962), .D(n4960), .S0(n5068), .S1(
        n5969), .Y(n4964) );
  MX4X2 U4596 ( .A(n4943), .B(n4941), .C(n4942), .D(n4940), .S0(n5068), .S1(
        n5969), .Y(n4944) );
  MX4X2 U4597 ( .A(n4958), .B(n4956), .C(n4957), .D(n4955), .S0(n5068), .S1(
        n5065), .Y(n4959) );
  MX4X2 U4598 ( .A(n4968), .B(n4966), .C(n4967), .D(n4965), .S0(n5068), .S1(
        n5969), .Y(n4969) );
  MX4X2 U4599 ( .A(n4973), .B(n4971), .C(n4972), .D(n4970), .S0(n5068), .S1(
        n5969), .Y(n4974) );
  AOI211XL U4600 ( .A0(n5935), .A1(n2941), .B0(n2950), .C0(n5887), .Y(n2949)
         );
  NAND2X4 U4601 ( .A(n5952), .B(n4675), .Y(n2939) );
  AOI211XL U4602 ( .A0(n5935), .A1(n3141), .B0(n3150), .C0(n5886), .Y(n3149)
         );
  NAND2X4 U4603 ( .A(n5954), .B(n4674), .Y(n3139) );
  OAI222X1 U4604 ( .A0(n6347), .A1(n5893), .B0(n3939), .B1(n3929), .C0(n697), 
        .C1(n3930), .Y(n4595) );
  AOI211XL U4605 ( .A0(n5935), .A1(n3931), .B0(n3940), .C0(n5889), .Y(n3939)
         );
  NAND2X8 U4606 ( .A(n5954), .B(n3930), .Y(n3929) );
  NAND2X8 U4607 ( .A(n5954), .B(n3535), .Y(n3534) );
  NAND2X8 U4608 ( .A(n5952), .B(n3574), .Y(n3573) );
  NAND2X8 U4609 ( .A(n5954), .B(n3613), .Y(n3612) );
  NAND2X8 U4610 ( .A(n5952), .B(n3774), .Y(n3773) );
  NAND2X8 U4611 ( .A(n5954), .B(n3813), .Y(n3812) );
  NAND2X8 U4612 ( .A(n5952), .B(n3891), .Y(n3890) );
  CLKINVX12 U4613 ( .A(n5670), .Y(n6353) );
  CLKINVX12 U4614 ( .A(n3930), .Y(n6347) );
  AOI211XL U4615 ( .A0(n5918), .A1(n6485), .B0(n1760), .C0(n5794), .Y(n1759)
         );
  CLKINVX12 U4616 ( .A(n1743), .Y(n6401) );
  NAND3X4 U4617 ( .A(n3980), .B(n4032), .C(n4033), .Y(n3981) );
  AND3X6 U4618 ( .A(N5342), .B(N5341), .C(N5343), .Y(n4033) );
  OAI31X4 U4619 ( .A0(n6193), .A1(n6192), .A2(n6191), .B0(n6190), .Y(N5341) );
  CLKBUFX2 U4620 ( .A(n5255), .Y(n5245) );
  NOR3BX1 U4621 ( .AN(n6219), .B(n6218), .C(n6203), .Y(n6204) );
  OAI222X4 U4622 ( .A0(n4011), .A1(n3975), .B0(n4012), .B1(n5668), .C0(n4000), 
        .C1(n166), .Y(n1007) );
  AOI221X4 U4623 ( .A0(n4667), .A1(n3982), .B0(n5929), .B1(n3983), .C0(n4014), 
        .Y(n4011) );
  BUFX16 U4624 ( .A(n1044), .Y(n4697) );
  NOR2BXL U4625 ( .AN(n3980), .B(n5668), .Y(n1044) );
  AOI221X1 U4626 ( .A0(n3594), .A1(n4701), .B0(n4697), .B1(n3605), .C0(n3606), 
        .Y(n3604) );
  AOI221X1 U4627 ( .A0(n3555), .A1(n4701), .B0(n4697), .B1(n3566), .C0(n3567), 
        .Y(n3565) );
  AOI221X1 U4628 ( .A0(n3633), .A1(n4701), .B0(n4697), .B1(n3644), .C0(n3645), 
        .Y(n3643) );
  OAI222X4 U4629 ( .A0(n4023), .A1(n3975), .B0(n4024), .B1(n5668), .C0(n4000), 
        .C1(n170), .Y(n4698) );
  OAI222X4 U4630 ( .A0(n4023), .A1(n3975), .B0(n4024), .B1(n5668), .C0(n4000), 
        .C1(n170), .Y(n1017) );
  OAI222X4 U4631 ( .A0(n4029), .A1(n3975), .B0(n4030), .B1(n5668), .C0(n4000), 
        .C1(n172), .Y(n1037) );
  NOR3BX2 U4632 ( .AN(n6093), .B(n6092), .C(n6077), .Y(n6078) );
  NOR3BX1 U4633 ( .AN(n6188), .B(n6187), .C(n6172), .Y(n6173) );
  OAI222X4 U4634 ( .A0(n4005), .A1(n3975), .B0(n4006), .B1(n5668), .C0(n4000), 
        .C1(n164), .Y(n1002) );
  AOI221XL U4635 ( .A0(N3355), .A1(n3982), .B0(n5935), .B1(n3983), .C0(n4008), 
        .Y(n4005) );
  NOR3BX1 U4636 ( .AN(n6125), .B(n6124), .C(n6109), .Y(n6110) );
  AOI211X2 U4637 ( .A0(n6108), .A1(n6120), .B0(n6107), .C0(n6123), .Y(n6109)
         );
  NAND2X4 U4638 ( .A(n5953), .B(n1743), .Y(n1742) );
  INVX3 U4639 ( .A(n1043), .Y(n4700) );
  CLKINVX20 U4640 ( .A(n4700), .Y(n4701) );
  OAI221X4 U4641 ( .A0(n5668), .A1(n3980), .B0(n3975), .B1(n5669), .C0(n5916), 
        .Y(n1043) );
  NOR3BX1 U4642 ( .AN(n6283), .B(n6282), .C(n6267), .Y(n6268) );
  AOI211X2 U4643 ( .A0(n6266), .A1(n6278), .B0(n6265), .C0(n6281), .Y(n6267)
         );
  NAND2X6 U4644 ( .A(n5952), .B(n3852), .Y(n3851) );
  OA21X2 U4645 ( .A0(n4053), .A1(n4696), .B0(n4036), .Y(n4825) );
  NOR2BX4 U4646 ( .AN(n5669), .B(n4036), .Y(n3982) );
  OR3X6 U4647 ( .A(n6112), .B(n6080), .C(n6144), .Y(n4036) );
  OAI22X1 U4648 ( .A0(n5913), .A1(n1854), .B0(n1866), .B1(n4637), .Y(n1865) );
  AOI221X4 U4649 ( .A0(n6598), .A1(n4696), .B0(n6533), .B1(n4650), .C0(n1691), 
        .Y(n1690) );
  AOI221X4 U4650 ( .A0(n6606), .A1(n4696), .B0(n6541), .B1(n4650), .C0(n1647), 
        .Y(n1646) );
  AOI221X4 U4651 ( .A0(n6590), .A1(n4696), .B0(n6525), .B1(n4650), .C0(n1735), 
        .Y(n1734) );
  OAI22X1 U4652 ( .A0(n5912), .A1(n3675), .B0(n3685), .B1(n4637), .Y(n3684) );
  OAI22X1 U4653 ( .A0(n976), .A1(n3758), .B0(n3768), .B1(n4637), .Y(n3767) );
  OAI22X1 U4654 ( .A0(n976), .A1(n3714), .B0(n3725), .B1(n4637), .Y(n3724) );
  OAI22X1 U4655 ( .A0(n5916), .A1(n3914), .B0(n3924), .B1(n4637), .Y(n3923) );
  OAI22X1 U4656 ( .A0(n5916), .A1(n3836), .B0(n3846), .B1(n4637), .Y(n3845) );
  OAI22X1 U4657 ( .A0(n976), .A1(n3797), .B0(n3807), .B1(n4637), .Y(n3806) );
  OAI22X1 U4658 ( .A0(n5916), .A1(n3875), .B0(n3885), .B1(n4637), .Y(n3884) );
  OAI22X1 U4659 ( .A0(n5913), .A1(n3597), .B0(n3607), .B1(n4637), .Y(n3606) );
  OAI22X1 U4660 ( .A0(n5915), .A1(n3558), .B0(n3568), .B1(n4637), .Y(n3567) );
  OAI22X1 U4661 ( .A0(n5914), .A1(n3636), .B0(n3646), .B1(n4637), .Y(n3645) );
  BUFX20 U4662 ( .A(n5447), .Y(n5448) );
  OAI22X1 U4663 ( .A0(n5916), .A1(n3953), .B0(n3964), .B1(n4637), .Y(n3963) );
  OAI22X1 U4664 ( .A0(n5913), .A1(n1765), .B0(n1779), .B1(n4637), .Y(n1778) );
  NAND2X2 U4665 ( .A(n1428), .B(n1432), .Y(n1080) );
  CLKBUFX3 U4666 ( .A(n1159), .Y(n4702) );
  CLKBUFX3 U4667 ( .A(n1108), .Y(n4703) );
  CLKBUFX3 U4668 ( .A(n1090), .Y(n4704) );
  NAND2X2 U4669 ( .A(n1428), .B(n1436), .Y(n1084) );
  CLKBUFX3 U4670 ( .A(n1155), .Y(n4705) );
  CLKBUFX3 U4671 ( .A(n1102), .Y(n4706) );
  CLKBUFX3 U4672 ( .A(n1082), .Y(n4707) );
  CLKBUFX3 U4673 ( .A(n1143), .Y(n4708) );
  NAND2X2 U4674 ( .A(n1475), .B(n1436), .Y(n1171) );
  NAND2X2 U4675 ( .A(n1433), .B(n1441), .Y(n1091) );
  CLKBUFX3 U4676 ( .A(n1116), .Y(n4709) );
  CLKBUFX3 U4677 ( .A(n1129), .Y(n4710) );
  CLKBUFX3 U4678 ( .A(n1157), .Y(n4711) );
  CLKBUFX3 U4679 ( .A(n1147), .Y(n4712) );
  NAND2X2 U4680 ( .A(n1475), .B(n1432), .Y(n1167) );
  CLKBUFX3 U4681 ( .A(n1118), .Y(n4713) );
  CLKBUFX3 U4682 ( .A(n1081), .Y(n4714) );
  NOR3X4 U4683 ( .A(n6691), .B(n6690), .C(n6692), .Y(n1435) );
  CLKBUFX3 U4684 ( .A(n1117), .Y(n4715) );
  CLKBUFX3 U4685 ( .A(n1141), .Y(n4716) );
  AND2X1 U4686 ( .A(n1435), .B(n1460), .Y(n1136) );
  INVX3 U4687 ( .A(n1136), .Y(n4717) );
  NAND2X2 U4688 ( .A(n1428), .B(n1433), .Y(n1083) );
  NOR3X4 U4689 ( .A(n6657), .B(n6688), .C(n6653), .Y(n1428) );
  CLKBUFX3 U4690 ( .A(n1156), .Y(n4718) );
  NAND2X2 U4691 ( .A(n1432), .B(n1441), .Y(n1094) );
  NAND2X1 U4692 ( .A(n1470), .B(n1436), .Y(n1159) );
  NAND2X2 U4693 ( .A(n1475), .B(n1434), .Y(n1169) );
  CLKBUFX3 U4694 ( .A(n1130), .Y(n4719) );
  AND2X1 U4695 ( .A(n1470), .B(n1433), .Y(n1158) );
  INVX3 U4696 ( .A(n1158), .Y(n4720) );
  AND2X1 U4697 ( .A(n1465), .B(n1435), .Y(n1148) );
  INVX3 U4698 ( .A(n1148), .Y(n4721) );
  NAND2X2 U4699 ( .A(n1475), .B(n1431), .Y(n1168) );
  NOR3X4 U4700 ( .A(n6657), .B(n6687), .C(n6658), .Y(n1475) );
  NAND2X1 U4701 ( .A(n1470), .B(n1432), .Y(n1155) );
  NAND2X2 U4702 ( .A(n1465), .B(n1429), .Y(n1142) );
  NOR3X4 U4703 ( .A(n6655), .B(n6692), .C(n6656), .Y(n1429) );
  AND2X1 U4704 ( .A(n1475), .B(n1433), .Y(n1170) );
  INVX3 U4705 ( .A(n1170), .Y(n4722) );
  NAND2X1 U4706 ( .A(n1428), .B(n1434), .Y(n1082) );
  NAND2X1 U4707 ( .A(n1451), .B(n1434), .Y(n1117) );
  NAND2X1 U4708 ( .A(n1434), .B(n1441), .Y(n1090) );
  NAND2X1 U4709 ( .A(n1470), .B(n1434), .Y(n1157) );
  NAND2X2 U4710 ( .A(n1434), .B(n1460), .Y(n1133) );
  NAND2X2 U4711 ( .A(n1465), .B(n1434), .Y(n1145) );
  NAND2X1 U4712 ( .A(n1451), .B(n1431), .Y(n1116) );
  NAND2X1 U4713 ( .A(n1428), .B(n1431), .Y(n1081) );
  NAND2X1 U4714 ( .A(n1470), .B(n1431), .Y(n1156) );
  NAND2X1 U4715 ( .A(n1446), .B(n1431), .Y(n1108) );
  NAND2X2 U4716 ( .A(n1431), .B(n1460), .Y(n1132) );
  NAND2X2 U4717 ( .A(n1465), .B(n1431), .Y(n1144) );
  NAND2X1 U4718 ( .A(n1460), .B(n1430), .Y(n1129) );
  NAND2X1 U4719 ( .A(n1429), .B(n1460), .Y(n1130) );
  NAND2X2 U4720 ( .A(n1433), .B(n1460), .Y(n1134) );
  INVX12 U4721 ( .A(n6664), .Y(IROM_A[4]) );
  INVX12 U4722 ( .A(n6661), .Y(IROM_A[1]) );
  INVX3 U4723 ( .A(n6676), .Y(n6661) );
  NAND2X1 U4724 ( .A(n1465), .B(n1436), .Y(n1147) );
  NAND2X1 U4725 ( .A(n1465), .B(n1432), .Y(n1143) );
  NAND2X1 U4726 ( .A(n1465), .B(n1430), .Y(n1141) );
  NAND2X2 U4727 ( .A(n1465), .B(n1433), .Y(n1146) );
  NAND2X1 U4728 ( .A(n1451), .B(n1433), .Y(n1118) );
  NAND2X1 U4729 ( .A(n1446), .B(n1433), .Y(n1102) );
  INVX12 U4730 ( .A(n6659), .Y(IROM_A[5]) );
  XOR2XL U4731 ( .A(\add_118/carry[5] ), .B(n6672), .Y(N3385) );
  INVX12 U4732 ( .A(n6662), .Y(IROM_A[2]) );
  INVX3 U4733 ( .A(n6675), .Y(n6662) );
  INVX12 U4734 ( .A(n6655), .Y(IRAM_A[1]) );
  NOR3X2 U4735 ( .A(n6654), .B(n6691), .C(n6656), .Y(n1432) );
  INVX12 U4736 ( .A(n6657), .Y(IRAM_A[3]) );
  INVX3 U4737 ( .A(n6689), .Y(n6657) );
  NOR3X2 U4738 ( .A(n6658), .B(n6689), .C(n6653), .Y(n1446) );
  BUFX12 U4739 ( .A(n6671), .Y(IROM_rd) );
  BUFX12 U4740 ( .A(n6680), .Y(IRAM_D[6]) );
  BUFX12 U4741 ( .A(n6679), .Y(IRAM_D[7]) );
  BUFX12 U4742 ( .A(n6681), .Y(IRAM_D[5]) );
  BUFX12 U4743 ( .A(n6682), .Y(IRAM_D[4]) );
  BUFX12 U4744 ( .A(n6683), .Y(IRAM_D[3]) );
  BUFX12 U4745 ( .A(n6684), .Y(IRAM_D[2]) );
  BUFX12 U4746 ( .A(n6685), .Y(IRAM_D[1]) );
  BUFX12 U4747 ( .A(n6686), .Y(IRAM_D[0]) );
  BUFX12 U4748 ( .A(n6678), .Y(IRAM_valid) );
  INVX12 U4749 ( .A(n6663), .Y(IROM_A[3]) );
  INVX12 U4750 ( .A(n6658), .Y(IRAM_A[4]) );
  NOR3X2 U4751 ( .A(n6689), .B(n6688), .C(n6653), .Y(n1451) );
  INVX12 U4752 ( .A(n6656), .Y(IRAM_A[2]) );
  NOR3X2 U4753 ( .A(n6654), .B(n6690), .C(n6655), .Y(n1434) );
  NOR3X2 U4754 ( .A(n6691), .B(n6690), .C(n6654), .Y(n1436) );
  INVX12 U4755 ( .A(n6653), .Y(IRAM_A[5]) );
  XOR2XL U4756 ( .A(\add_139/carry[5] ), .B(IRAM_A[5]), .Y(N3455) );
  NOR3X2 U4757 ( .A(n6689), .B(n6687), .C(n6658), .Y(n1470) );
  NOR3X2 U4758 ( .A(n6688), .B(n6687), .C(n6657), .Y(n1465) );
  NOR3X2 U4759 ( .A(n6688), .B(n6687), .C(n6689), .Y(n1460) );
  INVX12 U4760 ( .A(N3380), .Y(IROM_A[0]) );
  CLKINVX1 U4761 ( .A(n6677), .Y(N3380) );
  INVX12 U4762 ( .A(n6654), .Y(IRAM_A[0]) );
  NOR3X2 U4763 ( .A(n6692), .B(n6690), .C(n6655), .Y(n1433) );
  NOR3X2 U4764 ( .A(n6692), .B(n6691), .C(n6656), .Y(n1431) );
  OR2XL U4765 ( .A(n5669), .B(n5691), .Y(n4746) );
  OR2XL U4766 ( .A(n3986), .B(n5743), .Y(n4747) );
  NAND2X1 U4767 ( .A(n4746), .B(n4747), .Y(n4020) );
  NAND3BX4 U4768 ( .AN(n4035), .B(n5669), .C(n4036), .Y(n3986) );
  AOI221XL U4769 ( .A0(N3357), .A1(n3982), .B0(n5925), .B1(n3983), .C0(n4020), 
        .Y(n4017) );
  INVXL U4770 ( .A(N3324), .Y(n4748) );
  INVX3 U4771 ( .A(n4748), .Y(n4749) );
  NOR3BX2 U4772 ( .AN(n5673), .B(n6666), .C(n5270), .Y(n3732) );
  INVX3 U4773 ( .A(n6325), .Y(n6345) );
  OR2X1 U4774 ( .A(n6399), .B(n5858), .Y(n4750) );
  OR2X1 U4775 ( .A(n1848), .B(n1831), .Y(n4751) );
  OR2XL U4776 ( .A(n277), .B(n4643), .Y(n4752) );
  AOI211XL U4777 ( .A0(n5917), .A1(n6481), .B0(n1849), .C0(n5794), .Y(n1848)
         );
  OAI2BB1XL U4778 ( .A0N(N3323), .A1N(N3324), .B0(n5971), .Y(N3330) );
  OR2X1 U4779 ( .A(n6352), .B(n5857), .Y(n4754) );
  OR2X4 U4780 ( .A(n3752), .B(n3734), .Y(n4755) );
  OR2X1 U4781 ( .A(n661), .B(n3735), .Y(n4756) );
  NAND3X6 U4782 ( .A(n4754), .B(n4755), .C(n4756), .Y(n4559) );
  INVX12 U4783 ( .A(n3735), .Y(n6352) );
  OR2XL U4784 ( .A(n5780), .B(n3757), .Y(n4757) );
  OR2X1 U4785 ( .A(n4658), .B(n3770), .Y(n4758) );
  NAND3X1 U4786 ( .A(n4757), .B(n4758), .C(n3771), .Y(n3766) );
  AOI221X1 U4787 ( .A0(n3755), .A1(n4701), .B0(n4697), .B1(n3766), .C0(n3767), 
        .Y(n3765) );
  OR2X1 U4788 ( .A(n645), .B(n3652), .Y(n4761) );
  INVX12 U4789 ( .A(n3652), .Y(n6354) );
  NAND2X8 U4790 ( .A(n5952), .B(n3652), .Y(n3651) );
  CLKINVX12 U4791 ( .A(n4855), .Y(n3652) );
  NOR2X8 U4792 ( .A(n6416), .B(n4033), .Y(n1054) );
  AOI211X2 U4793 ( .A0(n6126), .A1(n6125), .B0(n6124), .C0(n6123), .Y(n6128)
         );
  OR2X1 U4794 ( .A(n6401), .B(n5894), .Y(n4764) );
  OR2X1 U4795 ( .A(n1751), .B(n1742), .Y(n4765) );
  OR2XL U4796 ( .A(n257), .B(n1743), .Y(n4766) );
  AOI211XL U4797 ( .A0(n5934), .A1(n6485), .B0(n1752), .C0(n5889), .Y(n1751)
         );
  CLKINVX12 U4798 ( .A(n4809), .Y(n1743) );
  BUFX8 U4799 ( .A(N3323), .Y(n5637) );
  NAND2X2 U4800 ( .A(n4770), .B(n6158), .Y(N5081) );
  CLKINVX1 U4801 ( .A(n6161), .Y(n4767) );
  CLKINVX1 U4802 ( .A(n6160), .Y(n4768) );
  CLKINVX1 U4803 ( .A(n6159), .Y(n4769) );
  NOR2X1 U4804 ( .A(n6163), .B(n5945), .Y(n6160) );
  CLKBUFX3 U4805 ( .A(n5444), .Y(n5451) );
  INVX6 U4806 ( .A(n5924), .Y(n5921) );
  NAND2X1 U4807 ( .A(n6510), .B(n4650), .Y(n4776) );
  NAND2X1 U4808 ( .A(n5945), .B(n6068), .Y(n6047) );
  INVX8 U4809 ( .A(n4807), .Y(n3968) );
  CLKBUFX3 U4810 ( .A(n5254), .Y(n5248) );
  CLKINVX12 U4811 ( .A(n4847), .Y(n2306) );
  CLKINVX12 U4812 ( .A(n4846), .Y(n2345) );
  CLKINVX12 U4813 ( .A(n4845), .Y(n2384) );
  CLKINVX12 U4814 ( .A(n4850), .Y(n2189) );
  CLKINVX12 U4815 ( .A(n4851), .Y(n2150) );
  CLKINVX12 U4816 ( .A(n4837), .Y(n2701) );
  CLKINVX12 U4817 ( .A(n4872), .Y(n2901) );
  CLKINVX12 U4818 ( .A(n4875), .Y(n2784) );
  CLKINVX12 U4819 ( .A(n4876), .Y(n2740) );
  INVX12 U4820 ( .A(n4881), .Y(n3813) );
  INVX12 U4821 ( .A(n4878), .Y(n3930) );
  INVX12 U4822 ( .A(n4879), .Y(n3891) );
  INVX12 U4823 ( .A(n4882), .Y(n3774) );
  INVX12 U4824 ( .A(n4880), .Y(n3852) );
  INVX12 U4825 ( .A(n4835), .Y(n1523) );
  INVX12 U4826 ( .A(n4836), .Y(n1479) );
  NAND2BX2 U4827 ( .AN(n5971), .B(n4771), .Y(n5973) );
  NOR2X1 U4828 ( .A(n5963), .B(n5955), .Y(n4771) );
  NAND3X1 U4829 ( .A(n4772), .B(n4773), .C(n4774), .Y(n4607) );
  OR2XL U4830 ( .A(n4027), .B(n3970), .Y(n4773) );
  BUFX4 U4831 ( .A(n5074), .Y(n5439) );
  AOI211X2 U4832 ( .A0(n6076), .A1(n6088), .B0(n6075), .C0(n6091), .Y(n6077)
         );
  NOR2X1 U4833 ( .A(n6068), .B(n5945), .Y(n6064) );
  OAI22X4 U4834 ( .A0(n5916), .A1(n4041), .B0(n4051), .B1(n4637), .Y(n4050) );
  CLKINVX6 U4835 ( .A(n1910), .Y(n6398) );
  CLKINVX1 U4836 ( .A(n4054), .Y(n6510) );
  OR2X1 U4837 ( .A(n6399), .B(n5864), .Y(n4777) );
  NOR2X2 U4838 ( .A(n1796), .B(n1787), .Y(n4784) );
  NOR2X2 U4839 ( .A(n6400), .B(n5895), .Y(n4783) );
  OR2XL U4840 ( .A(n3968), .B(n5858), .Y(n4772) );
  OR2XL U4841 ( .A(n709), .B(n6346), .Y(n4774) );
  NAND2XL U4842 ( .A(n6575), .B(n4696), .Y(n4775) );
  INVX1 U4843 ( .A(n6142), .Y(n6164) );
  OAI211XL U4844 ( .A0(N3358), .A1(n6083), .B0(n6082), .C0(n6081), .Y(n6085)
         );
  NAND2X4 U4845 ( .A(n5953), .B(n1871), .Y(n1870) );
  CLKBUFX4 U4846 ( .A(n5070), .Y(n5080) );
  NOR2BX1 U4847 ( .AN(n5941), .B(n5661), .Y(n6249) );
  NAND2BXL U4848 ( .AN(n5653), .B(n5659), .Y(n6093) );
  NAND2X8 U4849 ( .A(n5952), .B(n1910), .Y(n1909) );
  NAND3X1 U4850 ( .A(n4787), .B(n4788), .C(n4789), .Y(n4206) );
  AOI211XL U4851 ( .A0(n5920), .A1(n6473), .B0(n2003), .C0(n4698), .Y(n2002)
         );
  OR2XL U4852 ( .A(n2002), .B(n1987), .Y(n4788) );
  OR2XL U4853 ( .A(n276), .B(n4643), .Y(n4779) );
  AOI211XL U4854 ( .A0(n5920), .A1(n6481), .B0(n1847), .C0(n4698), .Y(n1846)
         );
  OR2X1 U4855 ( .A(n4832), .B(n5858), .Y(n4780) );
  OR2XL U4856 ( .A(n285), .B(n1871), .Y(n4782) );
  AOI211XL U4857 ( .A0(n5918), .A1(n6479), .B0(n1888), .C0(n5794), .Y(n1887)
         );
  CLKINVX12 U4858 ( .A(n4832), .Y(n1871) );
  NOR2XL U4859 ( .A(n265), .B(n1788), .Y(n4785) );
  OR3X2 U4860 ( .A(n4783), .B(n4784), .C(n4785), .Y(n4163) );
  AO21X4 U4861 ( .A0(n6094), .A1(n6093), .B0(n6092), .Y(n4786) );
  INVX1 U4862 ( .A(n6110), .Y(n6134) );
  NOR2X1 U4863 ( .A(n6165), .B(N3360), .Y(n6130) );
  NAND2X1 U4864 ( .A(n4667), .B(n4654), .Y(n6215) );
  INVX3 U4865 ( .A(n1988), .Y(n6396) );
  NAND2X1 U4866 ( .A(n5651), .B(n6101), .Y(n6095) );
  NOR2X1 U4867 ( .A(n6101), .B(n5651), .Y(n6097) );
  CLKINVX1 U4868 ( .A(n5673), .Y(n4822) );
  AND2X2 U4869 ( .A(n4892), .B(n4893), .Y(n4823) );
  NAND2X2 U4870 ( .A(n5954), .B(n1988), .Y(n1987) );
  NAND3X1 U4871 ( .A(n4793), .B(n4794), .C(n4795), .Y(n4191) );
  AOI211X1 U4872 ( .A0(n5917), .A1(n6477), .B0(n1927), .C0(n5794), .Y(n1926)
         );
  OR2X1 U4873 ( .A(n1926), .B(n1909), .Y(n4794) );
  MX4XL U4874 ( .A(n5018), .B(n5016), .C(n5017), .D(n5015), .S0(n5067), .S1(
        n5066), .Y(n5019) );
  MX4XL U4875 ( .A(\img_buff[60][6] ), .B(\img_buff[61][6] ), .C(
        \img_buff[62][6] ), .D(\img_buff[63][6] ), .S0(n5079), .S1(n5061), .Y(
        n5015) );
  MX4X4 U4876 ( .A(n5477), .B(n5475), .C(n5476), .D(n5474), .S0(n5649), .S1(
        n5269), .Y(n5478) );
  OR2X1 U4877 ( .A(n6396), .B(n5864), .Y(n4787) );
  OR2XL U4878 ( .A(n308), .B(n1988), .Y(n4789) );
  NAND2X2 U4879 ( .A(n4792), .B(n6095), .Y(N5079) );
  INVXL U4880 ( .A(n6097), .Y(n4790) );
  CLKINVX1 U4881 ( .A(n6096), .Y(n4791) );
  NAND3X6 U4882 ( .A(N5080), .B(N5079), .C(N5081), .Y(n4032) );
  CLKBUFX3 U4883 ( .A(n5776), .Y(n5779) );
  BUFX4 U4884 ( .A(n5443), .Y(n5453) );
  CLKBUFX2 U4885 ( .A(N3320), .Y(n5069) );
  NAND2X1 U4886 ( .A(n5948), .B(n6260), .Y(n6253) );
  INVX8 U4887 ( .A(n4806), .Y(n3980) );
  NOR2X1 U4888 ( .A(n6139), .B(n6150), .Y(n6151) );
  CLKBUFX3 U4889 ( .A(n6509), .Y(n5749) );
  NAND2X1 U4890 ( .A(n5658), .B(n6228), .Y(n6221) );
  NAND2X1 U4891 ( .A(n5651), .B(n6195), .Y(n6190) );
  OAI2BB1X1 U4892 ( .A0N(n6115), .A1N(N3358), .B0(n5665), .Y(n6114) );
  OAI2BB1XL U4893 ( .A0N(n6319), .A1N(n5665), .B0(n5922), .Y(n6241) );
  NOR2X1 U4894 ( .A(n6227), .B(N3353), .Y(n6223) );
  BUFX12 U4895 ( .A(n4673), .Y(n5958) );
  OAI2BB1XL U4896 ( .A0N(n6178), .A1N(n5665), .B0(n5657), .Y(n6177) );
  NOR2XL U4897 ( .A(n5946), .B(n5652), .Y(n6287) );
  NOR2XL U4898 ( .A(n6005), .B(N3353), .Y(n6001) );
  NAND2XL U4899 ( .A(N3360), .B(n6101), .Y(n6127) );
  INVX8 U4900 ( .A(n4841), .Y(n2545) );
  INVX8 U4901 ( .A(n4842), .Y(n2506) );
  INVX8 U4902 ( .A(n4843), .Y(n2467) );
  INVX8 U4903 ( .A(n4852), .Y(n2106) );
  INVX8 U4904 ( .A(n4839), .Y(n2623) );
  INVX8 U4905 ( .A(n4871), .Y(n2979) );
  INVX8 U4906 ( .A(n4870), .Y(n3018) );
  NAND2X4 U4907 ( .A(n5953), .B(n5670), .Y(n3690) );
  NOR2X8 U4908 ( .A(n93), .B(n6415), .Y(n978) );
  CLKBUFX3 U4909 ( .A(N3339), .Y(n5674) );
  OR2X1 U4910 ( .A(n6398), .B(n5858), .Y(n4793) );
  OR2XL U4911 ( .A(n293), .B(n1910), .Y(n4795) );
  INVXL U4912 ( .A(n6130), .Y(n4796) );
  CLKINVX1 U4913 ( .A(n6129), .Y(n4797) );
  NOR2X2 U4914 ( .A(n6170), .B(n6182), .Y(n6183) );
  AND3X2 U4915 ( .A(N4818), .B(N4817), .C(N4819), .Y(n4806) );
  NAND2BX2 U4916 ( .AN(n6287), .B(n6269), .Y(n6282) );
  NAND2X1 U4917 ( .A(n5929), .B(n6162), .Y(n6152) );
  INVX16 U4918 ( .A(n980), .Y(n6415) );
  NOR2X2 U4919 ( .A(n6258), .B(n5652), .Y(n6192) );
  OAI22X4 U4920 ( .A0(n3721), .A1(n4627), .B0(n1042), .B1(n3722), .Y(n3691) );
  BUFX20 U4921 ( .A(n3691), .Y(n5670) );
  OAI2BB1XL U4922 ( .A0N(n6209), .A1N(n5665), .B0(N3358), .Y(n6208) );
  NAND2BX1 U4923 ( .AN(n5926), .B(N3357), .Y(n6147) );
  NOR2BXL U4924 ( .AN(n5661), .B(n5941), .Y(n6337) );
  NAND3BX1 U4925 ( .AN(n5990), .B(n5989), .C(n5988), .Y(n5994) );
  NAND2BXL U4926 ( .AN(n5926), .B(n5656), .Y(n6264) );
  OAI2BB1X1 U4927 ( .A0N(n6083), .A1N(N3358), .B0(n5657), .Y(n6082) );
  NAND2BXL U4928 ( .AN(n5661), .B(n5941), .Y(n6339) );
  NOR2BX1 U4929 ( .AN(n5940), .B(n5659), .Y(n6154) );
  NOR2BXL U4930 ( .AN(n5653), .B(n5940), .Y(n6281) );
  BUFX8 U4931 ( .A(n5965), .Y(n5082) );
  CLKBUFX2 U4932 ( .A(n5965), .Y(n5442) );
  CLKBUFX4 U4933 ( .A(n5243), .Y(n5252) );
  CLKBUFX4 U4934 ( .A(n5269), .Y(n5267) );
  XNOR2XL U4935 ( .A(n5963), .B(\sub_80/carry[2] ), .Y(N3319) );
  MXI4X4 U4936 ( .A(n4914), .B(n4904), .C(n4909), .D(n4899), .S0(N3322), .S1(
        N3321), .Y(n4815) );
  INVX20 U4937 ( .A(n4818), .Y(N3322) );
  MX4X4 U4938 ( .A(n5582), .B(n5580), .C(n5581), .D(n5579), .S0(n5649), .S1(
        n5963), .Y(n5583) );
  AND2X2 U4939 ( .A(n978), .B(n989), .Y(n4802) );
  MX4XL U4940 ( .A(\img_buff[44][2] ), .B(\img_buff[45][2] ), .C(
        \img_buff[46][2] ), .D(\img_buff[47][2] ), .S0(n5441), .S1(n4632), .Y(
        n4940) );
  MX4XL U4941 ( .A(\img_buff[28][5] ), .B(\img_buff[29][5] ), .C(
        \img_buff[30][5] ), .D(\img_buff[31][5] ), .S0(n5078), .S1(n4631), .Y(
        n5005) );
  MX4XL U4942 ( .A(\img_buff[60][5] ), .B(\img_buff[61][5] ), .C(
        \img_buff[62][5] ), .D(\img_buff[63][5] ), .S0(n5078), .S1(n4695), .Y(
        n4995) );
  MX4XL U4943 ( .A(\img_buff[44][5] ), .B(\img_buff[45][5] ), .C(
        \img_buff[46][5] ), .D(\img_buff[47][5] ), .S0(n5250), .S1(n5262), .Y(
        n5188) );
  MX4XL U4944 ( .A(\img_buff[32][7] ), .B(\img_buff[33][7] ), .C(
        \img_buff[34][7] ), .D(\img_buff[35][7] ), .S0(n5081), .S1(n5056), .Y(
        n5043) );
  MX4XL U4945 ( .A(\img_buff[60][1] ), .B(\img_buff[61][1] ), .C(
        \img_buff[62][1] ), .D(\img_buff[63][1] ), .S0(n5434), .S1(n5443), .Y(
        n5293) );
  CLKBUFX3 U4946 ( .A(N3340), .Y(n5673) );
  CLKBUFX3 U4947 ( .A(N3340), .Y(n5672) );
  NOR3BX2 U4948 ( .AN(n5969), .B(n5966), .C(n5059), .Y(n1649) );
  NOR3BX2 U4949 ( .AN(n5959), .B(n5080), .C(n5960), .Y(n1650) );
  NOR3BX2 U4950 ( .AN(n5963), .B(n5966), .C(n4749), .Y(n1696) );
  NOR3BX2 U4951 ( .AN(n5963), .B(n5080), .C(n4749), .Y(n1695) );
  NOR3BX2 U4952 ( .AN(n5969), .B(n4636), .C(n5080), .Y(n1737) );
  NOR3BX2 U4953 ( .AN(n5963), .B(n5964), .C(n5966), .Y(n1784) );
  NOR3BX2 U4954 ( .AN(n5959), .B(n5961), .C(n5080), .Y(n1738) );
  NOR3BX2 U4955 ( .AN(n5963), .B(n5964), .C(n5080), .Y(n1785) );
  AND2X8 U4956 ( .A(n1053), .B(n4036), .Y(n1052) );
  OAI22XL U4957 ( .A0(n5669), .A1(n5679), .B0(n3986), .B1(n5730), .Y(n3995) );
  BUFX20 U4958 ( .A(n3985), .Y(n5669) );
  NAND3X6 U4959 ( .A(N3491), .B(N3490), .C(N3492), .Y(n3985) );
  AND2X2 U4960 ( .A(n5777), .B(n3980), .Y(n3978) );
  CLKBUFX3 U4961 ( .A(n5072), .Y(n5078) );
  CLKBUFX3 U4962 ( .A(n5072), .Y(n5077) );
  OA22X2 U4963 ( .A0(n1936), .A1(n5773), .B0(n5770), .B1(n1932), .Y(n1946) );
  OA22X2 U4964 ( .A0(n1814), .A1(n5773), .B0(n5770), .B1(n1810), .Y(n1825) );
  OA22X2 U4965 ( .A0(n1681), .A1(n4804), .B0(n5770), .B1(n1677), .Y(n1692) );
  OA22X2 U4966 ( .A0(n1725), .A1(n5772), .B0(n5770), .B1(n1721), .Y(n1736) );
  OA22X2 U4967 ( .A0(n1637), .A1(n5772), .B0(n5770), .B1(n1633), .Y(n1648) );
  NAND2X1 U4968 ( .A(n5930), .B(n6067), .Y(n6056) );
  OAI22X1 U4969 ( .A0(n5913), .A1(n1589), .B0(n1602), .B1(n4637), .Y(n1601) );
  OAI22X1 U4970 ( .A0(n5913), .A1(n1501), .B0(n1514), .B1(n4637), .Y(n1513) );
  OAI22X1 U4971 ( .A0(n5913), .A1(n1545), .B0(n1558), .B1(n4637), .Y(n1557) );
  NOR2X1 U4972 ( .A(n6075), .B(n6087), .Y(n6088) );
  CLKAND2X3 U4973 ( .A(n6074), .B(n6084), .Y(n6081) );
  NOR2X1 U4974 ( .A(n6070), .B(n5948), .Y(n6065) );
  AND2X2 U4975 ( .A(n6011), .B(n6021), .Y(n6018) );
  NAND2X1 U4976 ( .A(n5944), .B(n6163), .Y(n6143) );
  NOR2X1 U4977 ( .A(n6226), .B(n5655), .Y(n6181) );
  NOR2X1 U4978 ( .A(n6226), .B(n4667), .Y(n6212) );
  NAND2XL U4979 ( .A(N3364), .B(n5932), .Y(n6335) );
  OAI211XL U4980 ( .A0(n5657), .A1(n5987), .B0(n5986), .C0(n5985), .Y(n5989)
         );
  AOI31XL U4981 ( .A0(n5994), .A1(n5993), .A2(n5992), .B0(n5991), .Y(n5998) );
  NOR2X1 U4982 ( .A(n6228), .B(n5658), .Y(n6224) );
  NOR2X1 U4983 ( .A(n6195), .B(n5651), .Y(n6193) );
  NAND2XL U4984 ( .A(n6649), .B(n5669), .Y(n1048) );
  OAI2BB1XL U4985 ( .A0N(n6231), .A1N(n5922), .B0(n5665), .Y(n6329) );
  NOR2X1 U4986 ( .A(n6007), .B(n5658), .Y(n6002) );
  NOR2XL U4987 ( .A(n6070), .B(N3360), .Y(n6035) );
  OAI2BB1XL U4988 ( .A0N(n5987), .A1N(n5657), .B0(N3358), .Y(n5986) );
  INVX1 U4989 ( .A(N3333), .Y(n6574) );
  BUFX20 U4990 ( .A(N3366), .Y(n5665) );
  CLKBUFX3 U4991 ( .A(n5892), .Y(n5890) );
  BUFX20 U4992 ( .A(N3347), .Y(n5654) );
  OR2X2 U4993 ( .A(n5963), .B(\sub_80/carry[2] ), .Y(\sub_80/carry[3] ) );
  CLKAND2X6 U4994 ( .A(n6666), .B(n4894), .Y(n4820) );
  CLKXOR2X4 U4995 ( .A(n4819), .B(n5974), .Y(n4821) );
  MX4X1 U4996 ( .A(n5191), .B(n5189), .C(n5190), .D(n5188), .S0(n5271), .S1(
        n5268), .Y(n5192) );
  MX4X4 U4997 ( .A(n5206), .B(n5204), .C(n5205), .D(n5203), .S0(n5271), .S1(
        n5268), .Y(n5207) );
  MX4X1 U4998 ( .A(n5336), .B(n5334), .C(n5335), .D(n5333), .S0(n4800), .S1(
        n5959), .Y(n5337) );
  MX4XL U4999 ( .A(\img_buff[60][3] ), .B(\img_buff[61][3] ), .C(
        \img_buff[62][3] ), .D(\img_buff[63][3] ), .S0(n5435), .S1(n4699), .Y(
        n5333) );
  AOI211X1 U5000 ( .A0(N3375), .A1(n6497), .B0(n1496), .C0(n5794), .Y(n1495)
         );
  AOI211X1 U5001 ( .A0(n5926), .A1(n6497), .B0(n1492), .C0(n5869), .Y(n1491)
         );
  AOI211X1 U5002 ( .A0(n5929), .A1(n6497), .B0(n1490), .C0(n5879), .Y(n1489)
         );
  MX4X1 U5003 ( .A(\img_buff[32][3] ), .B(\img_buff[33][3] ), .C(
        \img_buff[34][3] ), .D(\img_buff[35][3] ), .S0(n5076), .S1(n5062), .Y(
        n4963) );
  MX4X1 U5004 ( .A(\img_buff[0][3] ), .B(\img_buff[1][3] ), .C(
        \img_buff[2][3] ), .D(\img_buff[3][3] ), .S0(n5434), .S1(n4699), .Y(
        n5351) );
  MX4XL U5005 ( .A(\img_buff[8][3] ), .B(\img_buff[9][3] ), .C(
        \img_buff[10][3] ), .D(\img_buff[11][3] ), .S0(n5076), .S1(n5063), .Y(
        n4971) );
  MX4X1 U5006 ( .A(n5116), .B(n5114), .C(n5115), .D(n5113), .S0(n5272), .S1(
        n5267), .Y(n5117) );
  MX4X1 U5007 ( .A(\img_buff[32][7] ), .B(\img_buff[33][7] ), .C(
        \img_buff[34][7] ), .D(\img_buff[35][7] ), .S0(n5440), .S1(n5454), .Y(
        n5421) );
  MX4XL U5008 ( .A(\img_buff[8][7] ), .B(\img_buff[9][7] ), .C(
        \img_buff[10][7] ), .D(\img_buff[11][7] ), .S0(n5081), .S1(n5063), .Y(
        n5051) );
  MX4XL U5009 ( .A(\img_buff[40][7] ), .B(\img_buff[41][7] ), .C(
        \img_buff[42][7] ), .D(\img_buff[43][7] ), .S0(n5081), .S1(n5062), .Y(
        n5041) );
  MX4X1 U5010 ( .A(\img_buff[0][3] ), .B(\img_buff[1][3] ), .C(
        \img_buff[2][3] ), .D(\img_buff[3][3] ), .S0(n5077), .S1(n5057), .Y(
        n4973) );
  MX4XL U5011 ( .A(\img_buff[0][3] ), .B(\img_buff[1][3] ), .C(
        \img_buff[2][3] ), .D(\img_buff[3][3] ), .S0(n5631), .S1(n5643), .Y(
        n5542) );
  MX4X1 U5012 ( .A(\img_buff[52][7] ), .B(\img_buff[53][7] ), .C(
        \img_buff[54][7] ), .D(\img_buff[55][7] ), .S0(n5252), .S1(n5264), .Y(
        n5225) );
  MX4X1 U5013 ( .A(\img_buff[32][7] ), .B(\img_buff[33][7] ), .C(
        \img_buff[34][7] ), .D(\img_buff[35][7] ), .S0(n5635), .S1(n5263), .Y(
        n5612) );
  MX4X1 U5014 ( .A(\img_buff[16][7] ), .B(\img_buff[17][7] ), .C(
        \img_buff[18][7] ), .D(\img_buff[19][7] ), .S0(n5635), .S1(n5263), .Y(
        n5617) );
  AND2XL U5015 ( .A(\img_buff[0][6] ), .B(n6415), .Y(n4801) );
  AND2XL U5016 ( .A(n4891), .B(n980), .Y(n4803) );
  INVX12 U5017 ( .A(n4828), .Y(n980) );
  BUFX20 U5018 ( .A(n1054), .Y(n5777) );
  CLKBUFX4 U5019 ( .A(n5627), .Y(n5628) );
  CLKBUFX4 U5020 ( .A(n5625), .Y(n5632) );
  NAND2BX2 U5021 ( .AN(n6255), .B(n6238), .Y(n6250) );
  OR3X4 U5022 ( .A(n6206), .B(n6175), .C(n6239), .Y(n4035) );
  CLKBUFX4 U5023 ( .A(n5072), .Y(n5074) );
  INVX3 U5024 ( .A(n5984), .Y(N3490) );
  INVX3 U5025 ( .A(n6048), .Y(N3492) );
  CLKBUFX4 U5026 ( .A(n5442), .Y(n5434) );
  CLKINVX1 U5027 ( .A(n3887), .Y(n6534) );
  CLKINVX1 U5028 ( .A(n3966), .Y(n6518) );
  CLKINVX1 U5029 ( .A(n3926), .Y(n6526) );
  CLKINVX1 U5030 ( .A(n3848), .Y(n6542) );
  CLKINVX1 U5031 ( .A(n3809), .Y(n6550) );
  CLKINVX1 U5032 ( .A(n3770), .Y(n6558) );
  CLKINVX1 U5033 ( .A(n3687), .Y(n6511) );
  INVX1 U5034 ( .A(n6268), .Y(n6289) );
  OAI22X1 U5035 ( .A0(n4639), .A1(n2329), .B0(n5785), .B1(n2335), .Y(n2340) );
  OAI22X1 U5036 ( .A0(n4638), .A1(n2251), .B0(n5785), .B1(n2257), .Y(n2262) );
  OAI22X1 U5037 ( .A0(n4639), .A1(n2368), .B0(n5785), .B1(n2374), .Y(n2379) );
  OAI22X1 U5038 ( .A0(n4640), .A1(n2407), .B0(n5785), .B1(n2413), .Y(n2418) );
  OAI22X1 U5039 ( .A0(n4638), .A1(n2446), .B0(n5785), .B1(n2452), .Y(n2458) );
  OAI22X1 U5040 ( .A0(n4639), .A1(n2290), .B0(n5785), .B1(n2296), .Y(n2301) );
  OAI22X1 U5041 ( .A0(n4639), .A1(n2212), .B0(n5785), .B1(n2218), .Y(n2223) );
  OAI22X1 U5042 ( .A0(n4640), .A1(n2173), .B0(n5785), .B1(n2179), .Y(n2184) );
  AOI221XL U5043 ( .A0(n6576), .A1(n4696), .B0(n6511), .B1(n4650), .C0(n3686), 
        .Y(n3685) );
  OAI22XL U5044 ( .A0(n5786), .A1(n3675), .B0(n5785), .B1(n3681), .Y(n3686) );
  OAI22XL U5045 ( .A0(n5786), .A1(n3758), .B0(n5782), .B1(n3764), .Y(n3769) );
  AOI221XL U5046 ( .A0(n6607), .A1(n4696), .B0(n6542), .B1(n4650), .C0(n3847), 
        .Y(n3846) );
  OAI22XL U5047 ( .A0(n5786), .A1(n3836), .B0(n5784), .B1(n3842), .Y(n3847) );
  AOI221XL U5048 ( .A0(n6615), .A1(n4696), .B0(n6550), .B1(n4650), .C0(n3808), 
        .Y(n3807) );
  OAI22XL U5049 ( .A0(n5786), .A1(n3797), .B0(n5784), .B1(n3803), .Y(n3808) );
  AOI221XL U5050 ( .A0(n6582), .A1(n4696), .B0(n6517), .B1(n4649), .C0(n1780), 
        .Y(n1779) );
  OAI22XL U5051 ( .A0(n5790), .A1(n1765), .B0(n5785), .B1(n1769), .Y(n1780) );
  OAI22XL U5052 ( .A0(n5790), .A1(n1677), .B0(n5785), .B1(n1681), .Y(n1691) );
  OAI22XL U5053 ( .A0(n5790), .A1(n1721), .B0(n5785), .B1(n1725), .Y(n1735) );
  OAI22XL U5054 ( .A0(n5790), .A1(n1633), .B0(n5785), .B1(n1637), .Y(n1647) );
  AOI221XL U5055 ( .A0(n6613), .A1(n4696), .B0(n6548), .B1(n4650), .C0(n1945), 
        .Y(n1944) );
  OAI22XL U5056 ( .A0(n5790), .A1(n1932), .B0(n5785), .B1(n1936), .Y(n1945) );
  OAI22XL U5057 ( .A0(n5790), .A1(n1893), .B0(n5785), .B1(n1897), .Y(n1906) );
  AOI221XL U5058 ( .A0(n6629), .A1(n4696), .B0(n6564), .B1(n4649), .C0(n1867), 
        .Y(n1866) );
  OAI22XL U5059 ( .A0(n5790), .A1(n1854), .B0(n5785), .B1(n1858), .Y(n1867) );
  AOI221XL U5060 ( .A0(n6637), .A1(n4696), .B0(n6572), .B1(n4649), .C0(n1824), 
        .Y(n1823) );
  OAI22XL U5061 ( .A0(n5790), .A1(n1810), .B0(n5785), .B1(n1814), .Y(n1824) );
  AOI221XL U5062 ( .A0(n6591), .A1(n4696), .B0(n6526), .B1(n4650), .C0(n3925), 
        .Y(n3924) );
  OAI22XL U5063 ( .A0(n5786), .A1(n3914), .B0(n5785), .B1(n3920), .Y(n3925) );
  AOI221XL U5064 ( .A0(n6583), .A1(n4696), .B0(n6518), .B1(n4650), .C0(n3965), 
        .Y(n3964) );
  OAI22XL U5065 ( .A0(n5786), .A1(n3953), .B0(n5785), .B1(n3959), .Y(n3965) );
  AOI221XL U5066 ( .A0(n6599), .A1(n4696), .B0(n6534), .B1(n4650), .C0(n3886), 
        .Y(n3885) );
  OAI22XL U5067 ( .A0(n5786), .A1(n3875), .B0(n5785), .B1(n3881), .Y(n3886) );
  INVX2 U5068 ( .A(n4814), .Y(n5755) );
  OAI221XL U5069 ( .A0(n5777), .A1(n1764), .B0(n4661), .B1(n1771), .C0(n1781), 
        .Y(n1777) );
  OAI221XL U5070 ( .A0(n5777), .A1(n1931), .B0(n4661), .B1(n1938), .C0(n1946), 
        .Y(n1942) );
  OAI221XL U5071 ( .A0(n5777), .A1(n1892), .B0(n4657), .B1(n1899), .C0(n1907), 
        .Y(n1903) );
  OAI221XL U5072 ( .A0(n5777), .A1(n1853), .B0(n4658), .B1(n1860), .C0(n1868), 
        .Y(n1864) );
  OAI221XL U5073 ( .A0(n5777), .A1(n1809), .B0(n4658), .B1(n1816), .C0(n1825), 
        .Y(n1821) );
  OAI221XL U5074 ( .A0(n5777), .A1(n2009), .B0(n4661), .B1(n2016), .C0(n2025), 
        .Y(n2021) );
  OAI221XL U5075 ( .A0(n5777), .A1(n1970), .B0(n4660), .B1(n1977), .C0(n1985), 
        .Y(n1981) );
  OAI221XL U5076 ( .A0(n5780), .A1(n3674), .B0(n4660), .B1(n3687), .C0(n3688), 
        .Y(n3683) );
  OA22XL U5077 ( .A0(n3681), .A1(n5773), .B0(n5768), .B1(n3675), .Y(n3688) );
  OA22XL U5078 ( .A0(n3764), .A1(n5773), .B0(n5769), .B1(n3758), .Y(n3771) );
  OAI221XL U5079 ( .A0(n5780), .A1(n3835), .B0(n4661), .B1(n3848), .C0(n3849), 
        .Y(n3844) );
  OA22XL U5080 ( .A0(n3842), .A1(n5773), .B0(n5771), .B1(n3836), .Y(n3849) );
  OAI221XL U5081 ( .A0(n5780), .A1(n3796), .B0(n4663), .B1(n3809), .C0(n3810), 
        .Y(n3805) );
  OA22XL U5082 ( .A0(n3803), .A1(n5773), .B0(n5771), .B1(n3797), .Y(n3810) );
  OAI221XL U5083 ( .A0(n5780), .A1(n3874), .B0(n4660), .B1(n3887), .C0(n3888), 
        .Y(n3883) );
  OA22XL U5084 ( .A0(n3881), .A1(n5772), .B0(n5771), .B1(n3875), .Y(n3888) );
  OA22XL U5085 ( .A0(n3603), .A1(n5772), .B0(n5767), .B1(n3597), .Y(n3610) );
  OA22XL U5086 ( .A0(n3642), .A1(n5772), .B0(n5769), .B1(n3636), .Y(n3649) );
  OA22XL U5087 ( .A0(n3564), .A1(n5772), .B0(n5767), .B1(n3558), .Y(n3571) );
  OAI221XL U5088 ( .A0(n5780), .A1(n3913), .B0(n4660), .B1(n3926), .C0(n3927), 
        .Y(n3922) );
  OA22XL U5089 ( .A0(n3920), .A1(n5772), .B0(n5771), .B1(n3914), .Y(n3927) );
  OAI221XL U5090 ( .A0(n5780), .A1(n3952), .B0(n4663), .B1(n3966), .C0(n3967), 
        .Y(n3962) );
  OA22XL U5091 ( .A0(n3959), .A1(n5772), .B0(n5771), .B1(n3953), .Y(n3967) );
  NOR2X2 U5092 ( .A(n6201), .B(n6213), .Y(n6214) );
  OAI22XL U5093 ( .A0(n5790), .A1(n1589), .B0(n5785), .B1(n1593), .Y(n1603) );
  AOI221XL U5094 ( .A0(n6630), .A1(n4696), .B0(n6565), .B1(n4650), .C0(n1515), 
        .Y(n1514) );
  OAI22XL U5095 ( .A0(n5790), .A1(n1501), .B0(n5785), .B1(n1505), .Y(n1515) );
  AOI221XL U5096 ( .A0(n6622), .A1(n4696), .B0(n6557), .B1(n4650), .C0(n1559), 
        .Y(n1558) );
  OAI22XL U5097 ( .A0(n5790), .A1(n1545), .B0(n5785), .B1(n1549), .Y(n1559) );
  OAI22XL U5098 ( .A0(n5786), .A1(n3519), .B0(n5785), .B1(n3525), .Y(n3530) );
  OAI22XL U5099 ( .A0(n5786), .A1(n3597), .B0(n5785), .B1(n3603), .Y(n3608) );
  OAI22XL U5100 ( .A0(n5786), .A1(n3636), .B0(n5785), .B1(n3642), .Y(n3647) );
  OAI22XL U5101 ( .A0(n5786), .A1(n3558), .B0(n5781), .B1(n3564), .Y(n3569) );
  AOI31X2 U5102 ( .A0(n6345), .A1(n6326), .A2(n6341), .B0(n6344), .Y(n6327) );
  NAND2BX2 U5103 ( .AN(n6129), .B(n6111), .Y(n6124) );
  NAND2BX2 U5104 ( .AN(n6223), .B(n6205), .Y(n6218) );
  NAND2BX2 U5105 ( .AN(n6192), .B(n6174), .Y(n6187) );
  AND2X2 U5106 ( .A(n6138), .B(n6147), .Y(n6145) );
  AND2X2 U5107 ( .A(n6321), .B(n6330), .Y(n6328) );
  INVX1 U5108 ( .A(n6173), .Y(n6196) );
  NOR3BX1 U5109 ( .AN(n6251), .B(n6250), .C(n6236), .Y(n6237) );
  OA22XL U5110 ( .A0(n3720), .A1(n5772), .B0(n5771), .B1(n3714), .Y(n3728) );
  INVX1 U5111 ( .A(n6296), .Y(n6317) );
  INVX1 U5112 ( .A(n5982), .Y(n6006) );
  NAND2BX2 U5113 ( .AN(n6096), .B(n6079), .Y(n6092) );
  OA22XL U5114 ( .A0(n1593), .A1(n5772), .B0(n5771), .B1(n1589), .Y(n1604) );
  OA22XL U5115 ( .A0(n1505), .A1(n5773), .B0(n5771), .B1(n1501), .Y(n1516) );
  OA22XL U5116 ( .A0(n1549), .A1(n5773), .B0(n5771), .B1(n1545), .Y(n1560) );
  INVX1 U5117 ( .A(n6015), .Y(n6038) );
  INVX3 U5118 ( .A(n6017), .Y(N3491) );
  CLKBUFX2 U5119 ( .A(N3323), .Y(n5636) );
  CLKBUFX2 U5120 ( .A(N3323), .Y(n5254) );
  NAND2XL U5121 ( .A(n5948), .B(n6070), .Y(n6062) );
  CLKINVX6 U5122 ( .A(n5932), .Y(n5928) );
  CLKBUFX2 U5123 ( .A(n5734), .Y(n5733) );
  NAND2X1 U5124 ( .A(n2461), .B(n1737), .Y(n2685) );
  NAND2X1 U5125 ( .A(n2144), .B(n1737), .Y(n2368) );
  NAND2X1 U5126 ( .A(n2144), .B(n1649), .Y(n2290) );
  NAND2X1 U5127 ( .A(n2461), .B(n1782), .Y(n2724) );
  NAND2X1 U5128 ( .A(n2461), .B(n1060), .Y(n2446) );
  NAND2X1 U5129 ( .A(n2144), .B(n1782), .Y(n2407) );
  NAND2X1 U5130 ( .A(n2144), .B(n1693), .Y(n2329) );
  NAND2X1 U5131 ( .A(n2144), .B(n1605), .Y(n2251) );
  NAND2X1 U5132 ( .A(n2144), .B(n1561), .Y(n2212) );
  NAND2X1 U5133 ( .A(n2144), .B(n1517), .Y(n2173) );
  NAND2X1 U5134 ( .A(n1826), .B(n1737), .Y(n2051) );
  NAND2X1 U5135 ( .A(n2461), .B(n1649), .Y(n2607) );
  NAND2X1 U5136 ( .A(n2461), .B(n1517), .Y(n2490) );
  NAND2X1 U5137 ( .A(n2461), .B(n1605), .Y(n2568) );
  NAND2X1 U5138 ( .A(n2461), .B(n1561), .Y(n2529) );
  NAND2X1 U5139 ( .A(n2144), .B(n1060), .Y(n2129) );
  NAND2X1 U5140 ( .A(n1826), .B(n1782), .Y(n2090) );
  NAND2X1 U5141 ( .A(n2461), .B(n1693), .Y(n2646) );
  NAND2X1 U5142 ( .A(n1059), .B(n1060), .Y(n1033) );
  NAND2X1 U5143 ( .A(n3729), .B(n1782), .Y(n4041) );
  NAND2X1 U5144 ( .A(n1061), .B(n1062), .Y(n1027) );
  NAND2X1 U5145 ( .A(n3729), .B(n1737), .Y(n3953) );
  NAND2X1 U5146 ( .A(n3095), .B(n1737), .Y(n3319) );
  NAND2X1 U5147 ( .A(n3729), .B(n1649), .Y(n3875) );
  NAND2X1 U5148 ( .A(n3095), .B(n1649), .Y(n3241) );
  NAND2X1 U5149 ( .A(n2778), .B(n1649), .Y(n2924) );
  NAND2X1 U5150 ( .A(n3729), .B(n1693), .Y(n3914) );
  NAND2X1 U5151 ( .A(n3729), .B(n1605), .Y(n3836) );
  NAND2X1 U5152 ( .A(n3729), .B(n1561), .Y(n3797) );
  NAND2X1 U5153 ( .A(n3729), .B(n1517), .Y(n3758) );
  NAND2X1 U5154 ( .A(n3412), .B(n1782), .Y(n3675) );
  NAND2X1 U5155 ( .A(n3412), .B(n1561), .Y(n3480) );
  NAND2X1 U5156 ( .A(n3412), .B(n1517), .Y(n3441) );
  NAND2X1 U5157 ( .A(n3412), .B(n1060), .Y(n3397) );
  NAND2X1 U5158 ( .A(n3095), .B(n1782), .Y(n3358) );
  NAND2X1 U5159 ( .A(n3095), .B(n1693), .Y(n3280) );
  NAND2X1 U5160 ( .A(n3095), .B(n1605), .Y(n3202) );
  NAND2X1 U5161 ( .A(n2778), .B(n1693), .Y(n2963) );
  NAND2X1 U5162 ( .A(n2778), .B(n1605), .Y(n2885) );
  NAND2X1 U5163 ( .A(n2778), .B(n1561), .Y(n2846) );
  NAND2X1 U5164 ( .A(n2778), .B(n1517), .Y(n2807) );
  NAND2X1 U5165 ( .A(n2778), .B(n1060), .Y(n2763) );
  NAND2X1 U5166 ( .A(n1826), .B(n1649), .Y(n1971) );
  NAND2X1 U5167 ( .A(n1826), .B(n1693), .Y(n2010) );
  INVX4 U5168 ( .A(n5835), .Y(n5831) );
  NAND2X1 U5169 ( .A(n3412), .B(n1737), .Y(n3636) );
  NAND2X1 U5170 ( .A(n2778), .B(n1737), .Y(n3002) );
  NAND2X1 U5171 ( .A(n3412), .B(n1649), .Y(n3558) );
  NAND2X1 U5172 ( .A(n3095), .B(n1517), .Y(n3124) );
  NAND2X1 U5173 ( .A(n3412), .B(n1605), .Y(n3519) );
  NAND2X1 U5174 ( .A(n3095), .B(n1561), .Y(n3163) );
  NAND2X1 U5175 ( .A(n3095), .B(n1060), .Y(n3080) );
  NAND2X1 U5176 ( .A(n2778), .B(n1782), .Y(n3041) );
  NAND2X1 U5177 ( .A(n3412), .B(n1693), .Y(n3597) );
  NAND2X1 U5178 ( .A(n1605), .B(n1059), .Y(n1589) );
  NAND2X1 U5179 ( .A(n1561), .B(n1059), .Y(n1545) );
  NAND2X1 U5180 ( .A(n1517), .B(n1059), .Y(n1501) );
  NAND2X1 U5181 ( .A(n3729), .B(n1060), .Y(n3714) );
  INVX3 U5182 ( .A(n5850), .Y(n5845) );
  INVX3 U5183 ( .A(n5822), .Y(n5819) );
  INVX3 U5184 ( .A(n5808), .Y(n5805) );
  INVX3 U5185 ( .A(n5798), .Y(n5806) );
  INVX3 U5186 ( .A(n5825), .Y(n5820) );
  INVX3 U5187 ( .A(n5824), .Y(n5821) );
  INVX3 U5188 ( .A(n5809), .Y(n5804) );
  INVX3 U5189 ( .A(n5810), .Y(n5800) );
  INVX3 U5190 ( .A(n5823), .Y(n5818) );
  INVX3 U5191 ( .A(n5849), .Y(n5847) );
  INVX3 U5192 ( .A(n5849), .Y(n5846) );
  INVX4 U5193 ( .A(n5828), .Y(n5834) );
  INVX4 U5194 ( .A(n5828), .Y(n5833) );
  INVX4 U5195 ( .A(n5828), .Y(n5832) );
  INVX3 U5196 ( .A(n5798), .Y(n5803) );
  INVX3 U5197 ( .A(n5798), .Y(n5802) );
  INVX3 U5198 ( .A(n5798), .Y(n5801) );
  INVX3 U5199 ( .A(n5798), .Y(n5799) );
  CLKINVX12 U5200 ( .A(n5956), .Y(n5955) );
  NAND3BXL U5201 ( .AN(n6086), .B(n6085), .C(n6084), .Y(n6090) );
  NAND2BX4 U5202 ( .AN(N3324), .B(n5965), .Y(n5971) );
  NAND2BXL U5203 ( .AN(n5656), .B(n5926), .Y(n6274) );
  AOI221X2 U5204 ( .A0(n3711), .A1(n4701), .B0(n4697), .B1(n3723), .C0(n3724), 
        .Y(n3721) );
  OAI2BB2X4 U5205 ( .B0(n4048), .B1(n4627), .A0N(n5667), .A1N(n971), .Y(n4807)
         );
  OA22X4 U5206 ( .A0(n1039), .A1(n4627), .B0(n1041), .B1(n1042), .Y(n4828) );
  NOR2BXL U5207 ( .AN(n5936), .B(n5654), .Y(n6043) );
  NOR2BXL U5208 ( .AN(n5457), .B(N3359), .Y(n6301) );
  NOR2BXL U5209 ( .AN(n5457), .B(N3351), .Y(n6273) );
  NOR2BXL U5210 ( .AN(n5654), .B(n5936), .Y(n6054) );
  NAND2BXL U5211 ( .AN(n5926), .B(N3357), .Y(n6293) );
  NAND2BXL U5212 ( .AN(n5940), .B(n5661), .Y(n6251) );
  NAND2BXL U5213 ( .AN(n5926), .B(n5656), .Y(n6051) );
  NAND2XL U5214 ( .A(n5655), .B(n5932), .Y(n6279) );
  AO21X2 U5215 ( .A0(n6036), .A1(n6009), .B0(n5665), .Y(n6008) );
  AOI31X2 U5216 ( .A0(n5993), .A1(n5978), .A2(n5977), .B0(n5990), .Y(n5980) );
  OAI211X2 U5217 ( .A0(n5976), .A1(n6003), .B0(n5975), .C0(n5985), .Y(n5977)
         );
  AO21X2 U5218 ( .A0(n6003), .A1(n5976), .B0(N3358), .Y(n5975) );
  NAND2BXL U5219 ( .AN(n5656), .B(n5926), .Y(n6042) );
  NAND2BXL U5220 ( .AN(n5653), .B(n5462), .Y(n6283) );
  NAND3BXL U5221 ( .AN(n6053), .B(n6052), .C(n6051), .Y(n6057) );
  OAI211XL U5222 ( .A0(n5657), .A1(n6262), .B0(n6050), .C0(n6049), .Y(n6052)
         );
  OAI2BB1XL U5223 ( .A0N(n4651), .A1N(N3358), .B0(n5922), .Y(n6146) );
  AND2XL U5224 ( .A(n5955), .B(\sub_80/carry[3] ), .Y(n4829) );
  NOR2BXL U5225 ( .AN(n5940), .B(n5653), .Y(n6058) );
  NOR2XL U5226 ( .A(n5949), .B(n5651), .Y(n6288) );
  NOR2XL U5227 ( .A(n5947), .B(N3353), .Y(n6315) );
  NAND2BXL U5228 ( .AN(n5941), .B(n5659), .Y(n6156) );
  NAND2XL U5229 ( .A(n4667), .B(n5932), .Y(n6307) );
  NAND2BXL U5230 ( .AN(n5940), .B(n5653), .Y(n6060) );
  NAND2BXL U5231 ( .AN(n5659), .B(n5941), .Y(n6311) );
  OAI2BB1XL U5232 ( .A0N(n6262), .A1N(n5657), .B0(n5922), .Y(n6050) );
  CLKBUFX2 U5233 ( .A(n5965), .Y(n5441) );
  NAND2XL U5234 ( .A(n5658), .B(n6007), .Y(n5999) );
  NAND2XL U5235 ( .A(n5658), .B(n5950), .Y(n6313) );
  NOR3X2 U5236 ( .A(N3333), .B(N3334), .C(n4800), .Y(n1061) );
  NOR3X2 U5237 ( .A(N3333), .B(N3334), .C(n5958), .Y(n1827) );
  NOR3X2 U5238 ( .A(n5958), .B(N3334), .C(n6574), .Y(n2462) );
  NOR3X2 U5239 ( .A(n4800), .B(N3334), .C(n6574), .Y(n2145) );
  NOR3X2 U5240 ( .A(N3327), .B(n4666), .C(n5270), .Y(n1063) );
  NOR3X2 U5241 ( .A(n5960), .B(n5959), .C(n5966), .Y(n1062) );
  NOR3X2 U5242 ( .A(n5634), .B(n5959), .C(n5961), .Y(n1606) );
  NOR3X2 U5243 ( .A(n5966), .B(n5959), .C(n5961), .Y(n1562) );
  NOR3X2 U5244 ( .A(n5960), .B(n5959), .C(n5634), .Y(n1518) );
  NAND2X1 U5245 ( .A(n3731), .B(n1739), .Y(n3959) );
  NAND2X1 U5246 ( .A(n3731), .B(n1695), .Y(n3920) );
  NAND2X1 U5247 ( .A(n3731), .B(n1651), .Y(n3881) );
  NAND2X1 U5248 ( .A(n3731), .B(n1607), .Y(n3842) );
  NAND2X1 U5249 ( .A(n3731), .B(n1563), .Y(n3803) );
  NAND2X1 U5250 ( .A(n3731), .B(n1519), .Y(n3764) );
  NAND2X1 U5251 ( .A(n3414), .B(n1784), .Y(n3681) );
  NAND2X1 U5252 ( .A(n3414), .B(n1563), .Y(n3486) );
  NAND2X1 U5253 ( .A(n3414), .B(n1519), .Y(n3447) );
  NAND2X1 U5254 ( .A(n3414), .B(n1064), .Y(n3403) );
  NAND2X1 U5255 ( .A(n3097), .B(n1784), .Y(n3364) );
  NAND2X1 U5256 ( .A(n3097), .B(n1739), .Y(n3325) );
  NAND2X1 U5257 ( .A(n3097), .B(n1695), .Y(n3286) );
  NAND2X1 U5258 ( .A(n3097), .B(n1651), .Y(n3247) );
  NAND2X1 U5259 ( .A(n3097), .B(n1607), .Y(n3208) );
  NAND2X1 U5260 ( .A(n2780), .B(n1695), .Y(n2969) );
  NAND2X1 U5261 ( .A(n2780), .B(n1651), .Y(n2930) );
  NAND2X1 U5262 ( .A(n2780), .B(n1607), .Y(n2891) );
  NAND2X1 U5263 ( .A(n2780), .B(n1563), .Y(n2852) );
  NAND2X1 U5264 ( .A(n2780), .B(n1519), .Y(n2813) );
  NAND2X1 U5265 ( .A(n2780), .B(n1064), .Y(n2769) );
  NAND2X1 U5266 ( .A(n3414), .B(n1739), .Y(n3642) );
  NAND2X1 U5267 ( .A(n3414), .B(n1695), .Y(n3603) );
  NAND2X1 U5268 ( .A(n3414), .B(n1651), .Y(n3564) );
  NAND2X1 U5269 ( .A(n3414), .B(n1607), .Y(n3525) );
  NAND2X1 U5270 ( .A(n3097), .B(n1563), .Y(n3169) );
  NAND2X1 U5271 ( .A(n3097), .B(n1519), .Y(n3130) );
  NAND2X1 U5272 ( .A(n3097), .B(n1064), .Y(n3086) );
  NAND2X1 U5273 ( .A(n2780), .B(n1784), .Y(n3047) );
  NAND2X1 U5274 ( .A(n2780), .B(n1739), .Y(n3008) );
  NAND2X1 U5275 ( .A(n3731), .B(n1784), .Y(n4047) );
  NAND2X1 U5276 ( .A(n3731), .B(n1064), .Y(n3720) );
  NAND2X1 U5277 ( .A(n1063), .B(n1064), .Y(n1032) );
  INVX1 U5278 ( .A(N3327), .Y(n6639) );
  NOR3X2 U5279 ( .A(N3327), .B(n4666), .C(n5955), .Y(n1828) );
  NOR3X2 U5280 ( .A(n5955), .B(n4666), .C(n6639), .Y(n2463) );
  NOR3X2 U5281 ( .A(n5270), .B(n4666), .C(n6639), .Y(n2146) );
  NAND2X1 U5282 ( .A(n1065), .B(n1066), .Y(n1025) );
  NAND2X1 U5283 ( .A(n1784), .B(n1063), .Y(n1769) );
  NAND2X1 U5284 ( .A(n1739), .B(n1063), .Y(n1725) );
  NAND2X1 U5285 ( .A(n1695), .B(n1063), .Y(n1681) );
  NAND2X1 U5286 ( .A(n1651), .B(n1063), .Y(n1637) );
  NAND2X1 U5287 ( .A(n1828), .B(n1064), .Y(n1814) );
  NAND2X1 U5288 ( .A(n1828), .B(n1563), .Y(n1897) );
  NAND2X1 U5289 ( .A(n1828), .B(n1607), .Y(n1936) );
  NAND2X1 U5290 ( .A(n1828), .B(n1519), .Y(n1858) );
  NAND2X1 U5291 ( .A(n1607), .B(n1063), .Y(n1593) );
  NAND2X1 U5292 ( .A(n1563), .B(n1063), .Y(n1549) );
  NAND2X1 U5293 ( .A(n1519), .B(n1063), .Y(n1505) );
  NAND2X1 U5294 ( .A(n1828), .B(n1695), .Y(n2014) );
  NAND2X1 U5295 ( .A(n1828), .B(n1651), .Y(n1975) );
  NAND2X1 U5296 ( .A(n2463), .B(n1784), .Y(n2730) );
  NAND2X1 U5297 ( .A(n2146), .B(n1784), .Y(n2413) );
  NAND2X1 U5298 ( .A(n2146), .B(n1695), .Y(n2335) );
  NAND2X1 U5299 ( .A(n2463), .B(n1064), .Y(n2452) );
  NAND2X1 U5300 ( .A(n2146), .B(n1563), .Y(n2218) );
  NAND2X1 U5301 ( .A(n2146), .B(n1607), .Y(n2257) );
  NAND2X1 U5302 ( .A(n2146), .B(n1519), .Y(n2179) );
  NAND2X1 U5303 ( .A(n2463), .B(n1739), .Y(n2691) );
  NAND2X1 U5304 ( .A(n2146), .B(n1739), .Y(n2374) );
  NAND2X1 U5305 ( .A(n2146), .B(n1651), .Y(n2296) );
  NAND2X1 U5306 ( .A(n1828), .B(n1784), .Y(n2096) );
  NAND2X1 U5307 ( .A(n2463), .B(n1695), .Y(n2652) );
  NAND2X1 U5308 ( .A(n2146), .B(n1064), .Y(n2135) );
  NAND2X1 U5309 ( .A(n2463), .B(n1563), .Y(n2535) );
  NAND2X1 U5310 ( .A(n2463), .B(n1607), .Y(n2574) );
  NAND2X1 U5311 ( .A(n2463), .B(n1519), .Y(n2496) );
  NAND2X1 U5312 ( .A(n1828), .B(n1739), .Y(n2057) );
  NAND2X1 U5313 ( .A(n2463), .B(n1651), .Y(n2613) );
  CLKINVX1 U5314 ( .A(n5818), .Y(n5826) );
  NAND2X1 U5315 ( .A(n1608), .B(n1065), .Y(n1588) );
  NAND2X1 U5316 ( .A(n1564), .B(n1065), .Y(n1544) );
  NAND2X1 U5317 ( .A(n1520), .B(n1065), .Y(n1500) );
  NAND2X1 U5318 ( .A(n1829), .B(n1696), .Y(n2009) );
  NAND2X1 U5319 ( .A(n1829), .B(n1066), .Y(n1809) );
  NAND2X1 U5320 ( .A(n1785), .B(n1065), .Y(n1764) );
  NAND2X1 U5321 ( .A(n1740), .B(n1065), .Y(n1720) );
  NAND2X1 U5322 ( .A(n1696), .B(n1065), .Y(n1676) );
  NAND2X1 U5323 ( .A(n1652), .B(n1065), .Y(n1632) );
  NAND2X1 U5324 ( .A(n1829), .B(n1564), .Y(n1892) );
  NAND2X1 U5325 ( .A(n1829), .B(n1608), .Y(n1931) );
  NAND2X1 U5326 ( .A(n1829), .B(n1520), .Y(n1853) );
  NAND2X1 U5327 ( .A(n1829), .B(n1652), .Y(n1970) );
  MXI4X4 U5328 ( .A(n5142), .B(n5132), .C(n5137), .D(n5127), .S0(n4666), .S1(
        N3327), .Y(n4808) );
  MX4X4 U5329 ( .A(n4954), .B(n4944), .C(n4949), .D(n4939), .S0(N3322), .S1(
        N3321), .Y(N3349) );
  MX4XL U5330 ( .A(n5361), .B(n5359), .C(n5360), .D(n5358), .S0(n4800), .S1(
        n5959), .Y(n5362) );
  MX4X4 U5331 ( .A(n5412), .B(n5402), .C(n5407), .D(n5397), .S0(N3334), .S1(
        N3333), .Y(N3361) );
  MX4XL U5332 ( .A(n5411), .B(n5409), .C(n5410), .D(n5408), .S0(n5957), .S1(
        n5456), .Y(n5412) );
  MX4XL U5333 ( .A(n5401), .B(n5399), .C(n5400), .D(n5398), .S0(n5957), .S1(
        n5456), .Y(n5402) );
  MX4XL U5334 ( .A(n5351), .B(n5349), .C(n5350), .D(n5348), .S0(n4800), .S1(
        n5959), .Y(n5352) );
  MX4XL U5335 ( .A(n5341), .B(n5339), .C(n5340), .D(n5338), .S0(n4800), .S1(
        n5959), .Y(n5342) );
  BUFX12 U5336 ( .A(N3350), .Y(n5657) );
  MX4XL U5337 ( .A(n4923), .B(n4921), .C(n4922), .D(n4920), .S0(n5067), .S1(
        n5065), .Y(n4924) );
  NAND2X8 U5338 ( .A(n5952), .B(n6346), .Y(n3970) );
  CLKINVX12 U5339 ( .A(n4867), .Y(n3179) );
  CLKINVX12 U5340 ( .A(n4865), .Y(n3257) );
  CLKINVX12 U5341 ( .A(n4864), .Y(n3296) );
  CLKINVX12 U5342 ( .A(n4863), .Y(n3335) );
  CLKINVX12 U5343 ( .A(n4860), .Y(n3457) );
  CLKINVX12 U5344 ( .A(n4861), .Y(n3418) );
  CLKINVX12 U5345 ( .A(n4862), .Y(n3374) );
  CLKINVX12 U5346 ( .A(n4866), .Y(n3218) );
  CLKINVX12 U5347 ( .A(n4854), .Y(n2028) );
  CLKINVX12 U5348 ( .A(n4853), .Y(n2067) );
  CLKINVX12 U5349 ( .A(n4868), .Y(n3101) );
  CLKINVX12 U5350 ( .A(n4869), .Y(n3057) );
  CLKINVX12 U5351 ( .A(n4859), .Y(n3496) );
  CLKINVX12 U5352 ( .A(n4830), .Y(n1949) );
  CLKINVX12 U5353 ( .A(n4857), .Y(n3574) );
  CLKINVX12 U5354 ( .A(n4856), .Y(n3613) );
  CLKINVX12 U5355 ( .A(n4858), .Y(n3535) );
  OA22X4 U5356 ( .A0(n1774), .A1(n4627), .B0(n1775), .B1(n1041), .Y(n4809) );
  OA22X4 U5357 ( .A0(n1686), .A1(n4627), .B0(n1041), .B1(n1687), .Y(n4810) );
  OA22X4 U5358 ( .A0(n1730), .A1(n4627), .B0(n1041), .B1(n1731), .Y(n4811) );
  OA22X4 U5359 ( .A0(n1642), .A1(n4627), .B0(n1041), .B1(n1643), .Y(n4812) );
  OA22X4 U5360 ( .A0(n2020), .A1(n4627), .B0(n1687), .B1(n1820), .Y(n4813) );
  OA22X4 U5361 ( .A0(n1598), .A1(n4627), .B0(n1041), .B1(n1599), .Y(n4834) );
  OA22X4 U5362 ( .A0(n1510), .A1(n4627), .B0(n1041), .B1(n1511), .Y(n4836) );
  OA22X4 U5363 ( .A0(n1554), .A1(n4627), .B0(n1041), .B1(n1555), .Y(n4835) );
  MX4X4 U5364 ( .A(n5312), .B(n5302), .C(n5307), .D(n5297), .S0(N3334), .S1(
        N3333), .Y(N3366) );
  MX4XL U5365 ( .A(n5301), .B(n5299), .C(n5300), .D(n5298), .S0(n5957), .S1(
        n5959), .Y(n5302) );
  MX4XL U5366 ( .A(n5296), .B(n5294), .C(n5295), .D(n5293), .S0(n5957), .S1(
        n5959), .Y(n5297) );
  MX4XL U5367 ( .A(n5391), .B(n5389), .C(n5390), .D(n5388), .S0(n4800), .S1(
        n5456), .Y(n5392) );
  MX4XL U5368 ( .A(n5381), .B(n5379), .C(n5380), .D(n5378), .S0(n4800), .S1(
        n5456), .Y(n5382) );
  MX4X4 U5369 ( .A(n4994), .B(n4984), .C(n4989), .D(n4979), .S0(N3322), .S1(
        N3321), .Y(N3347) );
  BUFX20 U5370 ( .A(N3367), .Y(n5666) );
  MX4XL U5371 ( .A(n5033), .B(n5031), .C(n5032), .D(n5030), .S0(n5067), .S1(
        n5066), .Y(n5034) );
  MX4XL U5372 ( .A(n5023), .B(n5021), .C(n5022), .D(n5020), .S0(n5067), .S1(
        n5066), .Y(n5024) );
  MX4XL U5373 ( .A(n5054), .B(n5044), .C(n5049), .D(n5039), .S0(N3322), .S1(
        N3321), .Y(N3344) );
  MX4XL U5374 ( .A(n5038), .B(n5036), .C(n5037), .D(n5035), .S0(n5069), .S1(
        n5066), .Y(n5039) );
  MX4XL U5375 ( .A(n5048), .B(n5046), .C(n5047), .D(n5045), .S0(n5068), .S1(
        n5066), .Y(n5049) );
  MX4X4 U5376 ( .A(n5432), .B(n5422), .C(n5427), .D(n5417), .S0(N3334), .S1(
        N3333), .Y(N3360) );
  MX4XL U5377 ( .A(n5416), .B(n5414), .C(n5415), .D(n5413), .S0(n4800), .S1(
        n5456), .Y(n5417) );
  MX4XL U5378 ( .A(n5426), .B(n5424), .C(n5425), .D(n5423), .S0(n5957), .S1(
        n5456), .Y(n5427) );
  XOR2X4 U5379 ( .A(n4819), .B(n4820), .Y(n4818) );
  CLKINVX12 U5380 ( .A(n4821), .Y(N3334) );
  MX4XL U5381 ( .A(n4998), .B(n4996), .C(n4997), .D(n4995), .S0(n5067), .S1(
        n5066), .Y(n4999) );
  MX4XL U5382 ( .A(n5008), .B(n5006), .C(n5007), .D(n5005), .S0(n5067), .S1(
        n5066), .Y(n5009) );
  MX4XL U5383 ( .A(n5607), .B(n5605), .C(n5606), .D(n5604), .S0(n5650), .S1(
        n5963), .Y(n5608) );
  AOI32XL U5384 ( .A0(n4064), .A1(n5964), .A2(n4066), .B0(n4749), .B1(n4067), 
        .Y(n4065) );
  OAI32XL U5385 ( .A0(n4085), .A1(n5955), .A2(reset), .B0(n4086), .B1(n5270), 
        .Y(n4612) );
  CLKINVX1 U5386 ( .A(n5815), .Y(n5827) );
  NAND3X2 U5387 ( .A(n6661), .B(n6662), .C(n6660), .Y(n1042) );
  OAI221XL U5388 ( .A0(n5635), .A1(n4073), .B0(n4068), .B1(n5438), .C0(n6648), 
        .Y(n4067) );
  NOR2XL U5389 ( .A(n5440), .B(n4073), .Y(n4069) );
  AOI211XL U5390 ( .A0(n5918), .A1(n3692), .B0(n3709), .C0(n4628), .Y(n3708)
         );
  AOI211XL U5391 ( .A0(n5925), .A1(n3692), .B0(n3705), .C0(n5866), .Y(n3704)
         );
  AOI211XL U5392 ( .A0(n5917), .A1(n3180), .B0(n3197), .C0(n4629), .Y(n3196)
         );
  AOI211XL U5393 ( .A0(n5917), .A1(n2941), .B0(n2958), .C0(n5792), .Y(n2957)
         );
  AOI211XL U5394 ( .A0(n5917), .A1(n2863), .B0(n2880), .C0(n5792), .Y(n2879)
         );
  AOI211XL U5395 ( .A0(n5926), .A1(n3180), .B0(n3193), .C0(n5866), .Y(n3192)
         );
  AOI211XL U5396 ( .A0(n5925), .A1(n2941), .B0(n2954), .C0(n5867), .Y(n2953)
         );
  AOI211XL U5397 ( .A0(n5926), .A1(n2863), .B0(n2876), .C0(n5867), .Y(n2875)
         );
  AOI211XL U5398 ( .A0(n5917), .A1(n2902), .B0(n2919), .C0(n5792), .Y(n2918)
         );
  AOI211XL U5399 ( .A0(n5917), .A1(n2824), .B0(n2841), .C0(n5792), .Y(n2840)
         );
  AOI211XL U5400 ( .A0(n5926), .A1(n2902), .B0(n2915), .C0(n5867), .Y(n2914)
         );
  AOI211XL U5401 ( .A0(n5926), .A1(n2824), .B0(n2837), .C0(n5867), .Y(n2836)
         );
  AOI211XL U5402 ( .A0(n5917), .A1(n3258), .B0(n3275), .C0(n4630), .Y(n3274)
         );
  AOI211XL U5403 ( .A0(n5926), .A1(n3258), .B0(n3271), .C0(n5867), .Y(n3270)
         );
  AOI211XL U5404 ( .A0(n5917), .A1(n3336), .B0(n3353), .C0(n4629), .Y(n3352)
         );
  AOI211XL U5405 ( .A0(n5917), .A1(n3297), .B0(n3314), .C0(n4630), .Y(n3313)
         );
  AOI211XL U5406 ( .A0(n5926), .A1(n3336), .B0(n3349), .C0(n5866), .Y(n3348)
         );
  AOI211XL U5407 ( .A0(n5926), .A1(n3297), .B0(n3310), .C0(n5867), .Y(n3309)
         );
  AOI211XL U5408 ( .A0(n5917), .A1(n3458), .B0(n3475), .C0(n4629), .Y(n3474)
         );
  AOI211XL U5409 ( .A0(n5917), .A1(n3419), .B0(n3436), .C0(n4630), .Y(n3435)
         );
  AOI211XL U5410 ( .A0(n5917), .A1(n3375), .B0(n3392), .C0(n4629), .Y(n3391)
         );
  AOI211XL U5411 ( .A0(n5917), .A1(n3219), .B0(n3236), .C0(n4630), .Y(n3235)
         );
  AOI211XL U5412 ( .A0(n5926), .A1(n3458), .B0(n3471), .C0(n5867), .Y(n3470)
         );
  AOI211XL U5413 ( .A0(n5926), .A1(n3419), .B0(n3432), .C0(n5866), .Y(n3431)
         );
  AOI211XL U5414 ( .A0(n5926), .A1(n3375), .B0(n3388), .C0(n5866), .Y(n3387)
         );
  AOI211XL U5415 ( .A0(n5926), .A1(n3219), .B0(n3232), .C0(n5867), .Y(n3231)
         );
  AOI211XL U5416 ( .A0(N3375), .A1(n3653), .B0(n3670), .C0(n5794), .Y(n3669)
         );
  AOI211XL U5417 ( .A0(n5926), .A1(n3653), .B0(n3666), .C0(n5866), .Y(n3665)
         );
  AOI211XL U5418 ( .A0(n5918), .A1(n3736), .B0(n3753), .C0(n4629), .Y(n3752)
         );
  AOI211XL U5419 ( .A0(n5926), .A1(n3736), .B0(n3749), .C0(n5866), .Y(n3748)
         );
  AOI211XL U5420 ( .A0(n5917), .A1(n3019), .B0(n3036), .C0(n4629), .Y(n3035)
         );
  AOI211XL U5421 ( .A0(n5917), .A1(n2980), .B0(n2997), .C0(n4630), .Y(n2996)
         );
  AOI211XL U5422 ( .A0(n5926), .A1(n3019), .B0(n3032), .C0(n5867), .Y(n3031)
         );
  AOI211XL U5423 ( .A0(n5926), .A1(n2980), .B0(n2993), .C0(n5866), .Y(n2992)
         );
  AOI211XL U5424 ( .A0(n5917), .A1(n3141), .B0(n3158), .C0(n4628), .Y(n3157)
         );
  AOI211XL U5425 ( .A0(n5917), .A1(n3102), .B0(n3119), .C0(n4629), .Y(n3118)
         );
  AOI211XL U5426 ( .A0(n5917), .A1(n3058), .B0(n3075), .C0(n4630), .Y(n3074)
         );
  AOI211XL U5427 ( .A0(n5925), .A1(n3141), .B0(n3154), .C0(n5866), .Y(n3153)
         );
  AOI211XL U5428 ( .A0(n5926), .A1(n3102), .B0(n3115), .C0(n5866), .Y(n3114)
         );
  AOI211XL U5429 ( .A0(n5926), .A1(n3058), .B0(n3071), .C0(n5867), .Y(n3070)
         );
  AOI211XL U5430 ( .A0(n5917), .A1(n3497), .B0(n3514), .C0(n4628), .Y(n3513)
         );
  AOI211XL U5431 ( .A0(n5926), .A1(n3497), .B0(n3510), .C0(n5866), .Y(n3509)
         );
  AOI211XL U5432 ( .A0(n5917), .A1(n3575), .B0(n3592), .C0(n4628), .Y(n3591)
         );
  AOI211XL U5433 ( .A0(n5926), .A1(n3575), .B0(n3588), .C0(n5866), .Y(n3587)
         );
  AOI211XL U5434 ( .A0(N3375), .A1(n3614), .B0(n3631), .C0(n4628), .Y(n3630)
         );
  AOI211XL U5435 ( .A0(n5459), .A1(n3614), .B0(n3627), .C0(n5866), .Y(n3626)
         );
  AOI211XL U5436 ( .A0(n5917), .A1(n3536), .B0(n3553), .C0(n5794), .Y(n3552)
         );
  AOI211XL U5437 ( .A0(n5459), .A1(n3536), .B0(n3549), .C0(n5866), .Y(n3548)
         );
  AOI211XL U5438 ( .A0(N3375), .A1(n3814), .B0(n3831), .C0(n4628), .Y(n3830)
         );
  AOI211XL U5439 ( .A0(n5459), .A1(n3814), .B0(n3827), .C0(n5866), .Y(n3826)
         );
  AOI211XL U5440 ( .A0(N3375), .A1(n3775), .B0(n3792), .C0(n4629), .Y(n3791)
         );
  AOI211XL U5441 ( .A0(n5459), .A1(n3775), .B0(n3788), .C0(n5866), .Y(n3787)
         );
  AOI211XL U5442 ( .A0(n5917), .A1(n3892), .B0(n3909), .C0(n5794), .Y(n3908)
         );
  AOI211XL U5443 ( .A0(n5459), .A1(n3892), .B0(n3905), .C0(n5866), .Y(n3904)
         );
  AOI211XL U5444 ( .A0(n5918), .A1(n3931), .B0(n3948), .C0(n4630), .Y(n3947)
         );
  AOI211XL U5445 ( .A0(n5926), .A1(n3931), .B0(n3944), .C0(n5866), .Y(n3943)
         );
  AOI211XL U5446 ( .A0(n5917), .A1(n3853), .B0(n3870), .C0(n5794), .Y(n3869)
         );
  AOI211XL U5447 ( .A0(n5926), .A1(n3853), .B0(n3866), .C0(n5866), .Y(n3865)
         );
  AOI211XL U5448 ( .A0(n5917), .A1(n3971), .B0(n4028), .C0(n5794), .Y(n4027)
         );
  AOI211XL U5449 ( .A0(n5926), .A1(n3971), .B0(n4016), .C0(n5866), .Y(n4015)
         );
  MX4XL U5450 ( .A(\img_buff[48][2] ), .B(\img_buff[49][2] ), .C(
        \img_buff[50][2] ), .D(\img_buff[51][2] ), .S0(n5966), .S1(n4762), .Y(
        n4938) );
  MX4XL U5451 ( .A(\img_buff[56][2] ), .B(\img_buff[57][2] ), .C(
        \img_buff[58][2] ), .D(\img_buff[59][2] ), .S0(n5434), .S1(n5063), .Y(
        n4936) );
  MX4XL U5452 ( .A(\img_buff[60][2] ), .B(\img_buff[61][2] ), .C(
        \img_buff[62][2] ), .D(\img_buff[63][2] ), .S0(n5070), .S1(n4762), .Y(
        n4935) );
  MX4XL U5453 ( .A(\img_buff[16][2] ), .B(\img_buff[17][2] ), .C(
        \img_buff[18][2] ), .D(\img_buff[19][2] ), .S0(n5075), .S1(n5061), .Y(
        n4948) );
  MX4XL U5454 ( .A(\img_buff[24][2] ), .B(\img_buff[25][2] ), .C(
        \img_buff[26][2] ), .D(\img_buff[27][2] ), .S0(n5075), .S1(n5970), .Y(
        n4946) );
  MX4XL U5455 ( .A(\img_buff[28][2] ), .B(\img_buff[29][2] ), .C(
        \img_buff[30][2] ), .D(\img_buff[31][2] ), .S0(n5075), .S1(n4762), .Y(
        n4945) );
  MX4XL U5456 ( .A(\img_buff[12][2] ), .B(\img_buff[13][2] ), .C(
        \img_buff[14][2] ), .D(\img_buff[15][2] ), .S0(n5075), .S1(n5062), .Y(
        n4950) );
  MX4XL U5457 ( .A(n5396), .B(n5394), .C(n5395), .D(n5393), .S0(n5957), .S1(
        n5456), .Y(n5397) );
  MX4XL U5458 ( .A(n5376), .B(n5374), .C(n5375), .D(n5373), .S0(n4800), .S1(
        n5456), .Y(n5377) );
  MX4XL U5459 ( .A(\img_buff[48][5] ), .B(\img_buff[49][5] ), .C(
        \img_buff[50][5] ), .D(\img_buff[51][5] ), .S0(n5437), .S1(n5451), .Y(
        n5376) );
  MX4XL U5460 ( .A(\img_buff[56][5] ), .B(\img_buff[57][5] ), .C(
        \img_buff[58][5] ), .D(\img_buff[59][5] ), .S0(n5437), .S1(n5451), .Y(
        n5374) );
  MX4XL U5461 ( .A(\img_buff[60][5] ), .B(\img_buff[61][5] ), .C(
        \img_buff[62][5] ), .D(\img_buff[63][5] ), .S0(n5437), .S1(n5451), .Y(
        n5373) );
  MX4XL U5462 ( .A(\img_buff[44][1] ), .B(\img_buff[45][1] ), .C(
        \img_buff[46][1] ), .D(\img_buff[47][1] ), .S0(n5434), .S1(n5450), .Y(
        n5298) );
  MX4XL U5463 ( .A(\img_buff[32][2] ), .B(\img_buff[33][2] ), .C(
        \img_buff[34][2] ), .D(\img_buff[35][2] ), .S0(n5075), .S1(n5060), .Y(
        n4943) );
  MX4XL U5464 ( .A(\img_buff[0][2] ), .B(\img_buff[1][2] ), .C(
        \img_buff[2][2] ), .D(\img_buff[3][2] ), .S0(n5075), .S1(n4632), .Y(
        n4953) );
  MX4XL U5465 ( .A(n5311), .B(n5309), .C(n5310), .D(n5308), .S0(n4800), .S1(
        n5959), .Y(n5312) );
  MX4XL U5466 ( .A(\img_buff[0][1] ), .B(\img_buff[1][1] ), .C(
        \img_buff[2][1] ), .D(\img_buff[3][1] ), .S0(n5435), .S1(n5448), .Y(
        n5311) );
  MX4XL U5467 ( .A(\img_buff[8][1] ), .B(\img_buff[9][1] ), .C(
        \img_buff[10][1] ), .D(\img_buff[11][1] ), .S0(n5435), .S1(n5448), .Y(
        n5309) );
  MX4XL U5468 ( .A(\img_buff[12][1] ), .B(\img_buff[13][1] ), .C(
        \img_buff[14][1] ), .D(\img_buff[15][1] ), .S0(n5435), .S1(n5448), .Y(
        n5308) );
  MX4XL U5469 ( .A(\img_buff[48][1] ), .B(\img_buff[49][1] ), .C(
        \img_buff[50][1] ), .D(\img_buff[51][1] ), .S0(n5434), .S1(n5450), .Y(
        n5296) );
  MX4XL U5470 ( .A(\img_buff[32][1] ), .B(\img_buff[33][1] ), .C(
        \img_buff[34][1] ), .D(\img_buff[35][1] ), .S0(n5434), .S1(n5450), .Y(
        n5301) );
  MX4XL U5471 ( .A(\img_buff[16][0] ), .B(\img_buff[17][0] ), .C(
        \img_buff[18][0] ), .D(\img_buff[19][0] ), .S0(n5628), .S1(n5640), .Y(
        n5477) );
  MX4XL U5472 ( .A(\img_buff[36][2] ), .B(\img_buff[37][2] ), .C(
        \img_buff[38][2] ), .D(\img_buff[39][2] ), .S0(n5075), .S1(n5057), .Y(
        n4942) );
  MX4XL U5473 ( .A(\img_buff[4][2] ), .B(\img_buff[5][2] ), .C(
        \img_buff[6][2] ), .D(\img_buff[7][2] ), .S0(n5075), .S1(n5062), .Y(
        n4952) );
  MX4XL U5474 ( .A(\img_buff[52][2] ), .B(\img_buff[53][2] ), .C(
        \img_buff[54][2] ), .D(\img_buff[55][2] ), .S0(n5070), .S1(n5064), .Y(
        n4937) );
  MX4XL U5475 ( .A(\img_buff[20][2] ), .B(\img_buff[21][2] ), .C(
        \img_buff[22][2] ), .D(\img_buff[23][2] ), .S0(n5075), .S1(n5060), .Y(
        n4947) );
  MX4XL U5476 ( .A(n5406), .B(n5404), .C(n5405), .D(n5403), .S0(n5957), .S1(
        n5456), .Y(n5407) );
  MX4XL U5477 ( .A(n5386), .B(n5384), .C(n5385), .D(n5383), .S0(n5957), .S1(
        n5456), .Y(n5387) );
  MX4XL U5478 ( .A(\img_buff[28][5] ), .B(\img_buff[29][5] ), .C(
        \img_buff[30][5] ), .D(\img_buff[31][5] ), .S0(n5437), .S1(n5451), .Y(
        n5383) );
  MX4XL U5479 ( .A(n5346), .B(n5344), .C(n5345), .D(n5343), .S0(n4800), .S1(
        n5959), .Y(n5347) );
  MX4XL U5480 ( .A(n5306), .B(n5304), .C(n5305), .D(n5303), .S0(n4800), .S1(
        n5959), .Y(n5307) );
  MX4XL U5481 ( .A(\img_buff[16][1] ), .B(\img_buff[17][1] ), .C(
        \img_buff[18][1] ), .D(\img_buff[19][1] ), .S0(n5435), .S1(n5448), .Y(
        n5306) );
  MX4XL U5482 ( .A(\img_buff[24][1] ), .B(\img_buff[25][1] ), .C(
        \img_buff[26][1] ), .D(\img_buff[27][1] ), .S0(n5435), .S1(n5448), .Y(
        n5304) );
  MX4XL U5483 ( .A(\img_buff[28][1] ), .B(\img_buff[29][1] ), .C(
        \img_buff[30][1] ), .D(\img_buff[31][1] ), .S0(n5435), .S1(n5448), .Y(
        n5303) );
  MX4XL U5484 ( .A(\img_buff[52][1] ), .B(\img_buff[53][1] ), .C(
        \img_buff[54][1] ), .D(\img_buff[55][1] ), .S0(n5434), .S1(n5443), .Y(
        n5295) );
  MX4XL U5485 ( .A(\img_buff[36][1] ), .B(\img_buff[37][1] ), .C(
        \img_buff[38][1] ), .D(\img_buff[39][1] ), .S0(n5434), .S1(n5450), .Y(
        n5300) );
  MX4XL U5486 ( .A(\img_buff[20][1] ), .B(\img_buff[21][1] ), .C(
        \img_buff[22][1] ), .D(\img_buff[23][1] ), .S0(n5435), .S1(n5448), .Y(
        n5305) );
  MX4XL U5487 ( .A(\img_buff[4][1] ), .B(\img_buff[5][1] ), .C(
        \img_buff[6][1] ), .D(\img_buff[7][1] ), .S0(n5435), .S1(n5448), .Y(
        n5310) );
  MX4XL U5488 ( .A(\img_buff[40][2] ), .B(\img_buff[41][2] ), .C(
        \img_buff[42][2] ), .D(\img_buff[43][2] ), .S0(n5075), .S1(n4631), .Y(
        n4941) );
  MX4XL U5489 ( .A(\img_buff[8][2] ), .B(\img_buff[9][2] ), .C(
        \img_buff[10][2] ), .D(\img_buff[11][2] ), .S0(n5075), .S1(n5058), .Y(
        n4951) );
  MX4XL U5490 ( .A(\img_buff[56][1] ), .B(\img_buff[57][1] ), .C(
        \img_buff[58][1] ), .D(\img_buff[59][1] ), .S0(n5434), .S1(n5443), .Y(
        n5294) );
  MX4XL U5491 ( .A(\img_buff[40][1] ), .B(\img_buff[41][1] ), .C(
        \img_buff[42][1] ), .D(\img_buff[43][1] ), .S0(n5434), .S1(n5450), .Y(
        n5299) );
  MX4XL U5492 ( .A(\img_buff[12][1] ), .B(\img_buff[13][1] ), .C(
        \img_buff[14][1] ), .D(\img_buff[15][1] ), .S0(n5250), .S1(n5641), .Y(
        n5499) );
  MX4XL U5493 ( .A(\img_buff[60][3] ), .B(\img_buff[61][3] ), .C(
        \img_buff[62][3] ), .D(\img_buff[63][3] ), .S0(n5629), .S1(n4749), .Y(
        n5524) );
  MX4XL U5494 ( .A(\img_buff[48][4] ), .B(\img_buff[49][4] ), .C(
        \img_buff[50][4] ), .D(\img_buff[51][4] ), .S0(n5631), .S1(n5643), .Y(
        n5547) );
  MX4XL U5495 ( .A(\img_buff[56][4] ), .B(\img_buff[57][4] ), .C(
        \img_buff[58][4] ), .D(\img_buff[59][4] ), .S0(n5631), .S1(n5643), .Y(
        n5545) );
  MX4XL U5496 ( .A(\img_buff[60][4] ), .B(\img_buff[61][4] ), .C(
        \img_buff[62][4] ), .D(\img_buff[63][4] ), .S0(n5631), .S1(n5643), .Y(
        n5544) );
  MX4XL U5497 ( .A(\img_buff[48][5] ), .B(\img_buff[49][5] ), .C(
        \img_buff[50][5] ), .D(\img_buff[51][5] ), .S0(n5632), .S1(n5644), .Y(
        n5567) );
  MX4XL U5498 ( .A(\img_buff[56][5] ), .B(\img_buff[57][5] ), .C(
        \img_buff[58][5] ), .D(\img_buff[59][5] ), .S0(n5632), .S1(n5644), .Y(
        n5565) );
  MX4XL U5499 ( .A(\img_buff[60][5] ), .B(\img_buff[61][5] ), .C(
        \img_buff[62][5] ), .D(\img_buff[63][5] ), .S0(n5632), .S1(n5644), .Y(
        n5564) );
  MX4XL U5500 ( .A(\img_buff[60][7] ), .B(\img_buff[61][7] ), .C(
        \img_buff[62][7] ), .D(\img_buff[63][7] ), .S0(n5439), .S1(n5453), .Y(
        n5413) );
  MX4XL U5501 ( .A(\img_buff[44][5] ), .B(\img_buff[45][5] ), .C(
        \img_buff[46][5] ), .D(\img_buff[47][5] ), .S0(n5437), .S1(n5451), .Y(
        n5378) );
  MX4XL U5502 ( .A(\img_buff[60][1] ), .B(\img_buff[61][1] ), .C(
        \img_buff[62][1] ), .D(\img_buff[63][1] ), .S0(n5074), .S1(n4632), .Y(
        n4915) );
  MX4XL U5503 ( .A(\img_buff[44][1] ), .B(\img_buff[45][1] ), .C(
        \img_buff[46][1] ), .D(\img_buff[47][1] ), .S0(n5074), .S1(n4695), .Y(
        n4920) );
  MX4XL U5504 ( .A(\img_buff[56][3] ), .B(\img_buff[57][3] ), .C(
        \img_buff[58][3] ), .D(\img_buff[59][3] ), .S0(n5250), .S1(n5259), .Y(
        n5144) );
  MX4XL U5505 ( .A(\img_buff[60][3] ), .B(\img_buff[61][3] ), .C(
        \img_buff[62][3] ), .D(\img_buff[63][3] ), .S0(n5250), .S1(n5259), .Y(
        n5143) );
  MX4XL U5506 ( .A(\img_buff[60][3] ), .B(\img_buff[61][3] ), .C(
        \img_buff[62][3] ), .D(\img_buff[63][3] ), .S0(n5075), .S1(n5970), .Y(
        n4955) );
  MX4XL U5507 ( .A(\img_buff[48][1] ), .B(\img_buff[49][1] ), .C(
        \img_buff[50][1] ), .D(\img_buff[51][1] ), .S0(n5248), .S1(n5257), .Y(
        n5106) );
  MX4XL U5508 ( .A(\img_buff[56][1] ), .B(\img_buff[57][1] ), .C(
        \img_buff[58][1] ), .D(\img_buff[59][1] ), .S0(n5248), .S1(n5257), .Y(
        n5104) );
  MX4XL U5509 ( .A(\img_buff[60][1] ), .B(\img_buff[61][1] ), .C(
        \img_buff[62][1] ), .D(\img_buff[63][1] ), .S0(n5248), .S1(n5257), .Y(
        n5103) );
  MX4XL U5510 ( .A(\img_buff[44][1] ), .B(\img_buff[45][1] ), .C(
        \img_buff[46][1] ), .D(\img_buff[47][1] ), .S0(n5248), .S1(n5257), .Y(
        n5108) );
  MX4XL U5511 ( .A(\img_buff[12][1] ), .B(\img_buff[13][1] ), .C(
        \img_buff[14][1] ), .D(\img_buff[15][1] ), .S0(n5249), .S1(n5258), .Y(
        n5118) );
  MX4XL U5512 ( .A(\img_buff[0][1] ), .B(\img_buff[1][1] ), .C(
        \img_buff[2][1] ), .D(\img_buff[3][1] ), .S0(n5629), .S1(n5641), .Y(
        n5502) );
  MX4XL U5513 ( .A(n5013), .B(n5011), .C(n5012), .D(n5010), .S0(n5067), .S1(
        n5066), .Y(n5014) );
  MX4XL U5514 ( .A(n5431), .B(n5429), .C(n5430), .D(n5428), .S0(n4800), .S1(
        n5456), .Y(n5432) );
  MX4XL U5515 ( .A(\img_buff[48][5] ), .B(\img_buff[49][5] ), .C(
        \img_buff[50][5] ), .D(\img_buff[51][5] ), .S0(n5078), .S1(n4762), .Y(
        n4998) );
  MX4XL U5516 ( .A(\img_buff[32][5] ), .B(\img_buff[33][5] ), .C(
        \img_buff[34][5] ), .D(\img_buff[35][5] ), .S0(n5437), .S1(n5451), .Y(
        n5381) );
  MX4XL U5517 ( .A(\img_buff[48][1] ), .B(\img_buff[49][1] ), .C(
        \img_buff[50][1] ), .D(\img_buff[51][1] ), .S0(n5074), .S1(n5064), .Y(
        n4918) );
  MX4XL U5518 ( .A(\img_buff[32][1] ), .B(\img_buff[33][1] ), .C(
        \img_buff[34][1] ), .D(\img_buff[35][1] ), .S0(n5074), .S1(n4695), .Y(
        n4923) );
  MX4XL U5519 ( .A(\img_buff[32][1] ), .B(\img_buff[33][1] ), .C(
        \img_buff[34][1] ), .D(\img_buff[35][1] ), .S0(n5248), .S1(n5257), .Y(
        n5111) );
  MX4XL U5520 ( .A(\img_buff[0][1] ), .B(\img_buff[1][1] ), .C(
        \img_buff[2][1] ), .D(\img_buff[3][1] ), .S0(n5249), .S1(n5258), .Y(
        n5121) );
  MX4XL U5521 ( .A(\img_buff[16][1] ), .B(\img_buff[17][1] ), .C(
        \img_buff[18][1] ), .D(\img_buff[19][1] ), .S0(n5436), .S1(n5063), .Y(
        n4928) );
  MX4XL U5522 ( .A(\img_buff[0][1] ), .B(\img_buff[1][1] ), .C(
        \img_buff[2][1] ), .D(\img_buff[3][1] ), .S0(n5436), .S1(n5057), .Y(
        n4933) );
  MX4XL U5523 ( .A(\img_buff[32][5] ), .B(\img_buff[33][5] ), .C(
        \img_buff[34][5] ), .D(\img_buff[35][5] ), .S0(n5078), .S1(n5970), .Y(
        n5003) );
  MX4XL U5524 ( .A(\img_buff[16][1] ), .B(\img_buff[17][1] ), .C(
        \img_buff[18][1] ), .D(\img_buff[19][1] ), .S0(n5626), .S1(n5641), .Y(
        n5497) );
  MX4XL U5525 ( .A(\img_buff[24][1] ), .B(\img_buff[25][1] ), .C(
        \img_buff[26][1] ), .D(\img_buff[27][1] ), .S0(n5244), .S1(n5641), .Y(
        n5495) );
  MX4XL U5526 ( .A(\img_buff[28][1] ), .B(\img_buff[29][1] ), .C(
        \img_buff[30][1] ), .D(\img_buff[31][1] ), .S0(n5624), .S1(n5641), .Y(
        n5494) );
  MX4XL U5527 ( .A(\img_buff[4][1] ), .B(\img_buff[5][1] ), .C(
        \img_buff[6][1] ), .D(\img_buff[7][1] ), .S0(n5250), .S1(n5641), .Y(
        n5501) );
  MX4XL U5528 ( .A(\img_buff[16][4] ), .B(\img_buff[17][4] ), .C(
        \img_buff[18][4] ), .D(\img_buff[19][4] ), .S0(n5631), .S1(n5643), .Y(
        n5557) );
  MX4XL U5529 ( .A(\img_buff[24][4] ), .B(\img_buff[25][4] ), .C(
        \img_buff[26][4] ), .D(\img_buff[27][4] ), .S0(n5631), .S1(n5643), .Y(
        n5555) );
  MX4XL U5530 ( .A(\img_buff[28][4] ), .B(\img_buff[29][4] ), .C(
        \img_buff[30][4] ), .D(\img_buff[31][4] ), .S0(n5631), .S1(n5643), .Y(
        n5554) );
  MX4XL U5531 ( .A(n5028), .B(n5026), .C(n5027), .D(n5025), .S0(n5067), .S1(
        n5066), .Y(n5029) );
  MX4XL U5532 ( .A(\img_buff[52][5] ), .B(\img_buff[53][5] ), .C(
        \img_buff[54][5] ), .D(\img_buff[55][5] ), .S0(n5078), .S1(n5061), .Y(
        n4997) );
  MX4XL U5533 ( .A(\img_buff[52][7] ), .B(\img_buff[53][7] ), .C(
        \img_buff[54][7] ), .D(\img_buff[55][7] ), .S0(n5439), .S1(n5453), .Y(
        n5415) );
  MX4XL U5534 ( .A(\img_buff[36][5] ), .B(\img_buff[37][5] ), .C(
        \img_buff[38][5] ), .D(\img_buff[39][5] ), .S0(n5437), .S1(n5451), .Y(
        n5380) );
  MX4XL U5535 ( .A(\img_buff[52][1] ), .B(\img_buff[53][1] ), .C(
        \img_buff[54][1] ), .D(\img_buff[55][1] ), .S0(n5074), .S1(n4631), .Y(
        n4917) );
  MX4XL U5536 ( .A(\img_buff[36][1] ), .B(\img_buff[37][1] ), .C(
        \img_buff[38][1] ), .D(\img_buff[39][1] ), .S0(n5074), .S1(n5055), .Y(
        n4922) );
  MX4XL U5537 ( .A(\img_buff[36][5] ), .B(\img_buff[37][5] ), .C(
        \img_buff[38][5] ), .D(\img_buff[39][5] ), .S0(n5247), .S1(n5262), .Y(
        n5190) );
  MX4XL U5538 ( .A(\img_buff[16][1] ), .B(\img_buff[17][1] ), .C(
        \img_buff[18][1] ), .D(\img_buff[19][1] ), .S0(n5249), .S1(n5258), .Y(
        n5116) );
  MX4XL U5539 ( .A(\img_buff[24][1] ), .B(\img_buff[25][1] ), .C(
        \img_buff[26][1] ), .D(\img_buff[27][1] ), .S0(n5249), .S1(n5258), .Y(
        n5114) );
  MX4XL U5540 ( .A(\img_buff[28][1] ), .B(\img_buff[29][1] ), .C(
        \img_buff[30][1] ), .D(\img_buff[31][1] ), .S0(n5249), .S1(n5258), .Y(
        n5113) );
  MX4XL U5541 ( .A(\img_buff[36][1] ), .B(\img_buff[37][1] ), .C(
        \img_buff[38][1] ), .D(\img_buff[39][1] ), .S0(n5248), .S1(n5257), .Y(
        n5110) );
  MX4XL U5542 ( .A(\img_buff[4][1] ), .B(\img_buff[5][1] ), .C(
        \img_buff[6][1] ), .D(\img_buff[7][1] ), .S0(n5249), .S1(n5258), .Y(
        n5120) );
  MX4XL U5543 ( .A(\img_buff[52][5] ), .B(\img_buff[53][5] ), .C(
        \img_buff[54][5] ), .D(\img_buff[55][5] ), .S0(n5437), .S1(n5451), .Y(
        n5375) );
  MX4XL U5544 ( .A(\img_buff[20][1] ), .B(\img_buff[21][1] ), .C(
        \img_buff[22][1] ), .D(\img_buff[23][1] ), .S0(n5626), .S1(n5641), .Y(
        n5496) );
  MX4XL U5545 ( .A(\img_buff[52][1] ), .B(\img_buff[53][1] ), .C(
        \img_buff[54][1] ), .D(\img_buff[55][1] ), .S0(n5628), .S1(n5640), .Y(
        n5486) );
  MX4XL U5546 ( .A(\img_buff[36][1] ), .B(\img_buff[37][1] ), .C(
        \img_buff[38][1] ), .D(\img_buff[39][1] ), .S0(n5628), .S1(n5640), .Y(
        n5491) );
  MX4XL U5547 ( .A(\img_buff[52][4] ), .B(\img_buff[53][4] ), .C(
        \img_buff[54][4] ), .D(\img_buff[55][4] ), .S0(n5631), .S1(n5643), .Y(
        n5546) );
  MX4XL U5548 ( .A(\img_buff[20][4] ), .B(\img_buff[21][4] ), .C(
        \img_buff[22][4] ), .D(\img_buff[23][4] ), .S0(n5631), .S1(n5643), .Y(
        n5556) );
  MX4XL U5549 ( .A(\img_buff[36][4] ), .B(\img_buff[37][4] ), .C(
        \img_buff[38][4] ), .D(\img_buff[39][4] ), .S0(n5631), .S1(n5643), .Y(
        n5551) );
  MX4XL U5550 ( .A(\img_buff[52][1] ), .B(\img_buff[53][1] ), .C(
        \img_buff[54][1] ), .D(\img_buff[55][1] ), .S0(n5248), .S1(n5257), .Y(
        n5105) );
  MX4XL U5551 ( .A(\img_buff[20][1] ), .B(\img_buff[21][1] ), .C(
        \img_buff[22][1] ), .D(\img_buff[23][1] ), .S0(n5249), .S1(n5258), .Y(
        n5115) );
  MX4XL U5552 ( .A(\img_buff[52][5] ), .B(\img_buff[53][5] ), .C(
        \img_buff[54][5] ), .D(\img_buff[55][5] ), .S0(n5632), .S1(n5644), .Y(
        n5566) );
  MX4XL U5553 ( .A(\img_buff[36][5] ), .B(\img_buff[37][5] ), .C(
        \img_buff[38][5] ), .D(\img_buff[39][5] ), .S0(n5632), .S1(n5644), .Y(
        n5571) );
  MX4XL U5554 ( .A(\img_buff[52][5] ), .B(\img_buff[53][5] ), .C(
        \img_buff[54][5] ), .D(\img_buff[55][5] ), .S0(n5244), .S1(n5262), .Y(
        n5185) );
  MX4XL U5555 ( .A(\img_buff[8][1] ), .B(\img_buff[9][1] ), .C(
        \img_buff[10][1] ), .D(\img_buff[11][1] ), .S0(n5250), .S1(n5641), .Y(
        n5500) );
  MX4XL U5556 ( .A(\img_buff[56][3] ), .B(\img_buff[57][3] ), .C(
        \img_buff[58][3] ), .D(\img_buff[59][3] ), .S0(n5637), .S1(n4749), .Y(
        n5525) );
  MX4XL U5557 ( .A(\img_buff[32][4] ), .B(\img_buff[33][4] ), .C(
        \img_buff[34][4] ), .D(\img_buff[35][4] ), .S0(n5631), .S1(n5643), .Y(
        n5552) );
  MX4XL U5558 ( .A(\img_buff[40][4] ), .B(\img_buff[41][4] ), .C(
        \img_buff[42][4] ), .D(\img_buff[43][4] ), .S0(n5631), .S1(n5643), .Y(
        n5550) );
  MX4XL U5559 ( .A(\img_buff[44][4] ), .B(\img_buff[45][4] ), .C(
        \img_buff[46][4] ), .D(\img_buff[47][4] ), .S0(n5631), .S1(n5643), .Y(
        n5549) );
  MX4X2 U5560 ( .A(n5572), .B(n5570), .C(n5571), .D(n5569), .S0(n5650), .S1(
        n5963), .Y(n5573) );
  MX4XL U5561 ( .A(\img_buff[32][5] ), .B(\img_buff[33][5] ), .C(
        \img_buff[34][5] ), .D(\img_buff[35][5] ), .S0(n5632), .S1(n5644), .Y(
        n5572) );
  MX4XL U5562 ( .A(\img_buff[40][5] ), .B(\img_buff[41][5] ), .C(
        \img_buff[42][5] ), .D(\img_buff[43][5] ), .S0(n5632), .S1(n5644), .Y(
        n5570) );
  MX4XL U5563 ( .A(\img_buff[44][5] ), .B(\img_buff[45][5] ), .C(
        \img_buff[46][5] ), .D(\img_buff[47][5] ), .S0(n5632), .S1(n5644), .Y(
        n5569) );
  MX4XL U5564 ( .A(n5003), .B(n5001), .C(n5002), .D(n5000), .S0(n5067), .S1(
        n5066), .Y(n5004) );
  MX4XL U5565 ( .A(\img_buff[44][5] ), .B(\img_buff[45][5] ), .C(
        \img_buff[46][5] ), .D(\img_buff[47][5] ), .S0(n5078), .S1(n5063), .Y(
        n5000) );
  MX4XL U5566 ( .A(\img_buff[36][5] ), .B(\img_buff[37][5] ), .C(
        \img_buff[38][5] ), .D(\img_buff[39][5] ), .S0(n5078), .S1(n5970), .Y(
        n5002) );
  MX4XL U5567 ( .A(\img_buff[40][5] ), .B(\img_buff[41][5] ), .C(
        \img_buff[42][5] ), .D(\img_buff[43][5] ), .S0(n5078), .S1(n5055), .Y(
        n5001) );
  MX4XL U5568 ( .A(n5421), .B(n5419), .C(n5420), .D(n5418), .S0(n4800), .S1(
        n5456), .Y(n5422) );
  MX4XL U5569 ( .A(\img_buff[56][5] ), .B(\img_buff[57][5] ), .C(
        \img_buff[58][5] ), .D(\img_buff[59][5] ), .S0(n5078), .S1(n5063), .Y(
        n4996) );
  MX4XL U5570 ( .A(\img_buff[56][7] ), .B(\img_buff[57][7] ), .C(
        \img_buff[58][7] ), .D(\img_buff[59][7] ), .S0(n5439), .S1(n5453), .Y(
        n5414) );
  MX4XL U5571 ( .A(\img_buff[40][5] ), .B(\img_buff[41][5] ), .C(
        \img_buff[42][5] ), .D(\img_buff[43][5] ), .S0(n5437), .S1(n5451), .Y(
        n5379) );
  MX4XL U5572 ( .A(\img_buff[56][1] ), .B(\img_buff[57][1] ), .C(
        \img_buff[58][1] ), .D(\img_buff[59][1] ), .S0(n5074), .S1(n5056), .Y(
        n4916) );
  MX4XL U5573 ( .A(\img_buff[40][1] ), .B(\img_buff[41][1] ), .C(
        \img_buff[42][1] ), .D(\img_buff[43][1] ), .S0(n5074), .S1(n5056), .Y(
        n4921) );
  MX4XL U5574 ( .A(\img_buff[40][5] ), .B(\img_buff[41][5] ), .C(
        \img_buff[42][5] ), .D(\img_buff[43][5] ), .S0(n5250), .S1(n5262), .Y(
        n5189) );
  MX4XL U5575 ( .A(\img_buff[56][3] ), .B(\img_buff[57][3] ), .C(
        \img_buff[58][3] ), .D(\img_buff[59][3] ), .S0(n5075), .S1(n5057), .Y(
        n4956) );
  MX4XL U5576 ( .A(\img_buff[40][1] ), .B(\img_buff[41][1] ), .C(
        \img_buff[42][1] ), .D(\img_buff[43][1] ), .S0(n5248), .S1(n5257), .Y(
        n5109) );
  MX4XL U5577 ( .A(\img_buff[8][1] ), .B(\img_buff[9][1] ), .C(
        \img_buff[10][1] ), .D(\img_buff[11][1] ), .S0(n5249), .S1(n5258), .Y(
        n5119) );
  MX4XL U5578 ( .A(\img_buff[48][1] ), .B(\img_buff[49][1] ), .C(
        \img_buff[50][1] ), .D(\img_buff[51][1] ), .S0(n5628), .S1(n5640), .Y(
        n5487) );
  MX4XL U5579 ( .A(\img_buff[56][1] ), .B(\img_buff[57][1] ), .C(
        \img_buff[58][1] ), .D(\img_buff[59][1] ), .S0(n5628), .S1(n5640), .Y(
        n5485) );
  MX4XL U5580 ( .A(\img_buff[60][1] ), .B(\img_buff[61][1] ), .C(
        \img_buff[62][1] ), .D(\img_buff[63][1] ), .S0(n5628), .S1(n5640), .Y(
        n5484) );
  MX4XL U5581 ( .A(\img_buff[32][1] ), .B(\img_buff[33][1] ), .C(
        \img_buff[34][1] ), .D(\img_buff[35][1] ), .S0(n5628), .S1(n5640), .Y(
        n5492) );
  MX4XL U5582 ( .A(\img_buff[40][1] ), .B(\img_buff[41][1] ), .C(
        \img_buff[42][1] ), .D(\img_buff[43][1] ), .S0(n5628), .S1(n5640), .Y(
        n5490) );
  MX4XL U5583 ( .A(\img_buff[44][1] ), .B(\img_buff[45][1] ), .C(
        \img_buff[46][1] ), .D(\img_buff[47][1] ), .S0(n5628), .S1(n5640), .Y(
        n5489) );
  MX4XL U5584 ( .A(\img_buff[60][7] ), .B(\img_buff[61][7] ), .C(
        \img_buff[62][7] ), .D(\img_buff[63][7] ), .S0(n5634), .S1(n5646), .Y(
        n5604) );
  MX4XL U5585 ( .A(\img_buff[60][7] ), .B(\img_buff[61][7] ), .C(
        \img_buff[62][7] ), .D(\img_buff[63][7] ), .S0(n5080), .S1(n5058), .Y(
        n5035) );
  MX4XL U5586 ( .A(n5622), .B(n5620), .C(n5621), .D(n5619), .S0(n5650), .S1(
        n5963), .Y(n5623) );
  MX4XL U5587 ( .A(n5053), .B(n5051), .C(n5052), .D(n5050), .S0(N3320), .S1(
        n5066), .Y(n5054) );
  MX4XL U5588 ( .A(\img_buff[32][5] ), .B(\img_buff[33][5] ), .C(
        \img_buff[34][5] ), .D(\img_buff[35][5] ), .S0(n5250), .S1(n5262), .Y(
        n5191) );
  MX4XL U5589 ( .A(n5617), .B(n5615), .C(n5616), .D(n5614), .S0(n5649), .S1(
        n5963), .Y(n5618) );
  MX4XL U5590 ( .A(\img_buff[52][7] ), .B(\img_buff[53][7] ), .C(
        \img_buff[54][7] ), .D(\img_buff[55][7] ), .S0(n5634), .S1(n5646), .Y(
        n5606) );
  MX4XL U5591 ( .A(\img_buff[52][7] ), .B(\img_buff[53][7] ), .C(
        \img_buff[54][7] ), .D(\img_buff[55][7] ), .S0(n5080), .S1(n4762), .Y(
        n5037) );
  MX4XL U5592 ( .A(n5612), .B(n5610), .C(n5611), .D(n5609), .S0(n5650), .S1(
        n5963), .Y(n5613) );
  MX4XL U5593 ( .A(\img_buff[56][7] ), .B(\img_buff[57][7] ), .C(
        \img_buff[58][7] ), .D(\img_buff[59][7] ), .S0(n5634), .S1(n5646), .Y(
        n5605) );
  MX4XL U5594 ( .A(n5043), .B(n5041), .C(n5042), .D(n5040), .S0(N3320), .S1(
        n5066), .Y(n5044) );
  MX4XL U5595 ( .A(\img_buff[56][7] ), .B(\img_buff[57][7] ), .C(
        \img_buff[58][7] ), .D(\img_buff[59][7] ), .S0(n5080), .S1(n4695), .Y(
        n5036) );
  NOR2X1 U5596 ( .A(n963), .B(cmd_reg[2]), .Y(n4058) );
  NAND3X1 U5597 ( .A(n4057), .B(n964), .C(cmd_reg[3]), .Y(n1028) );
  NAND3X1 U5598 ( .A(cmd_reg[3]), .B(n964), .C(n4058), .Y(n1035) );
  OAI21X1 U5599 ( .A0(n975), .A1(n93), .B0(n6642), .Y(n4064) );
  NOR2X1 U5600 ( .A(n964), .B(cmd_reg[3]), .Y(n4059) );
  NAND3X1 U5601 ( .A(cmd_reg[3]), .B(cmd_reg[0]), .C(n4058), .Y(n1031) );
  INVX1 U5602 ( .A(n6677), .Y(n6660) );
  NAND3X2 U5603 ( .A(n4059), .B(n963), .C(cmd_reg[2]), .Y(n3975) );
  OAI22XL U5604 ( .A0(n4712), .A1(n285), .B0(n4721), .B1(n277), .Y(n1461) );
  OAI22XL U5605 ( .A0(n4702), .A1(n349), .B0(n1160), .B1(n341), .Y(n1466) );
  OAI22XL U5606 ( .A0(n4712), .A1(n284), .B0(n4721), .B1(n276), .Y(n1407) );
  OAI22XL U5607 ( .A0(n4702), .A1(n348), .B0(n1160), .B1(n340), .Y(n1411) );
  OAI22XL U5608 ( .A0(n4712), .A1(n283), .B0(n4721), .B1(n275), .Y(n1366) );
  OAI22XL U5609 ( .A0(n4702), .A1(n347), .B0(n1160), .B1(n339), .Y(n1370) );
  OAI22XL U5610 ( .A0(n4712), .A1(n282), .B0(n4721), .B1(n274), .Y(n1325) );
  OAI22XL U5611 ( .A0(n4702), .A1(n346), .B0(n1160), .B1(n338), .Y(n1329) );
  OAI22XL U5612 ( .A0(n4712), .A1(n281), .B0(n4721), .B1(n273), .Y(n1284) );
  OAI22XL U5613 ( .A0(n4702), .A1(n345), .B0(n1160), .B1(n337), .Y(n1288) );
  OAI22XL U5614 ( .A0(n4712), .A1(n280), .B0(n4721), .B1(n272), .Y(n1243) );
  OAI22XL U5615 ( .A0(n4702), .A1(n344), .B0(n1160), .B1(n336), .Y(n1247) );
  OAI22XL U5616 ( .A0(n4712), .A1(n278), .B0(n4721), .B1(n270), .Y(n1137) );
  OAI22XL U5617 ( .A0(n4702), .A1(n342), .B0(n1160), .B1(n334), .Y(n1149) );
  OAI22XL U5618 ( .A0(n4712), .A1(n279), .B0(n4721), .B1(n271), .Y(n1202) );
  OAI22XL U5619 ( .A0(n4702), .A1(n343), .B0(n1160), .B1(n335), .Y(n1206) );
  OAI22XL U5620 ( .A0(n1171), .A1(n413), .B0(n1172), .B1(n405), .Y(n1471) );
  OAI22XL U5621 ( .A0(n1171), .A1(n412), .B0(n1172), .B1(n404), .Y(n1415) );
  OAI22XL U5622 ( .A0(n1171), .A1(n411), .B0(n1172), .B1(n403), .Y(n1374) );
  OAI22XL U5623 ( .A0(n1171), .A1(n410), .B0(n1172), .B1(n402), .Y(n1333) );
  OAI22XL U5624 ( .A0(n1171), .A1(n409), .B0(n1172), .B1(n401), .Y(n1292) );
  OAI22XL U5625 ( .A0(n1171), .A1(n408), .B0(n1172), .B1(n400), .Y(n1251) );
  OAI22XL U5626 ( .A0(n1171), .A1(n406), .B0(n1172), .B1(n398), .Y(n1161) );
  OAI22XL U5627 ( .A0(n1171), .A1(n407), .B0(n1172), .B1(n399), .Y(n1210) );
  OAI22XL U5628 ( .A0(n1084), .A1(n541), .B0(n1085), .B1(n533), .Y(n1424) );
  OAI22XL U5629 ( .A0(n1084), .A1(n540), .B0(n1085), .B1(n532), .Y(n1383) );
  OAI22XL U5630 ( .A0(n1084), .A1(n539), .B0(n1085), .B1(n531), .Y(n1342) );
  OAI22XL U5631 ( .A0(n1084), .A1(n538), .B0(n1085), .B1(n530), .Y(n1301) );
  OAI22XL U5632 ( .A0(n1084), .A1(n537), .B0(n1085), .B1(n529), .Y(n1260) );
  OAI22XL U5633 ( .A0(n1084), .A1(n536), .B0(n1085), .B1(n528), .Y(n1219) );
  OAI22XL U5634 ( .A0(n1084), .A1(n534), .B0(n1085), .B1(n526), .Y(n1074) );
  OAI22XL U5635 ( .A0(n1084), .A1(n535), .B0(n1085), .B1(n527), .Y(n1178) );
  OAI22XL U5636 ( .A0(n4708), .A1(n317), .B0(n1144), .B1(n309), .Y(n1463) );
  OAI22XL U5637 ( .A0(n4705), .A1(n381), .B0(n4718), .B1(n373), .Y(n1468) );
  OAI22XL U5638 ( .A0(n4708), .A1(n316), .B0(n1144), .B1(n308), .Y(n1409) );
  OAI22XL U5639 ( .A0(n4705), .A1(n380), .B0(n4718), .B1(n372), .Y(n1413) );
  OAI22XL U5640 ( .A0(n4708), .A1(n315), .B0(n1144), .B1(n307), .Y(n1368) );
  OAI22XL U5641 ( .A0(n4705), .A1(n379), .B0(n4718), .B1(n371), .Y(n1372) );
  OAI22XL U5642 ( .A0(n4708), .A1(n314), .B0(n1144), .B1(n306), .Y(n1327) );
  OAI22XL U5643 ( .A0(n4705), .A1(n378), .B0(n4718), .B1(n370), .Y(n1331) );
  OAI22XL U5644 ( .A0(n4708), .A1(n313), .B0(n1144), .B1(n305), .Y(n1286) );
  OAI22XL U5645 ( .A0(n4705), .A1(n377), .B0(n4718), .B1(n369), .Y(n1290) );
  OAI22XL U5646 ( .A0(n4708), .A1(n312), .B0(n1144), .B1(n304), .Y(n1245) );
  OAI22XL U5647 ( .A0(n4705), .A1(n376), .B0(n4718), .B1(n368), .Y(n1249) );
  OAI22XL U5648 ( .A0(n4708), .A1(n310), .B0(n1144), .B1(n302), .Y(n1139) );
  OAI22XL U5649 ( .A0(n4705), .A1(n374), .B0(n4718), .B1(n366), .Y(n1151) );
  OAI22XL U5650 ( .A0(n4708), .A1(n311), .B0(n1144), .B1(n303), .Y(n1204) );
  OAI22XL U5651 ( .A0(n4705), .A1(n375), .B0(n4718), .B1(n367), .Y(n1208) );
  OAI22XL U5652 ( .A0(n1145), .A1(n301), .B0(n1146), .B1(n293), .Y(n1462) );
  OAI22XL U5653 ( .A0(n4711), .A1(n365), .B0(n4720), .B1(n357), .Y(n1467) );
  OAI22XL U5654 ( .A0(n1145), .A1(n300), .B0(n1146), .B1(n292), .Y(n1408) );
  OAI22XL U5655 ( .A0(n4711), .A1(n364), .B0(n4720), .B1(n356), .Y(n1412) );
  OAI22XL U5656 ( .A0(n1145), .A1(n299), .B0(n1146), .B1(n291), .Y(n1367) );
  OAI22XL U5657 ( .A0(n4711), .A1(n363), .B0(n4720), .B1(n355), .Y(n1371) );
  OAI22XL U5658 ( .A0(n1145), .A1(n298), .B0(n1146), .B1(n290), .Y(n1326) );
  OAI22XL U5659 ( .A0(n4711), .A1(n362), .B0(n4720), .B1(n354), .Y(n1330) );
  OAI22XL U5660 ( .A0(n1145), .A1(n297), .B0(n1146), .B1(n289), .Y(n1285) );
  OAI22XL U5661 ( .A0(n4711), .A1(n361), .B0(n4720), .B1(n353), .Y(n1289) );
  OAI22XL U5662 ( .A0(n1145), .A1(n296), .B0(n1146), .B1(n288), .Y(n1244) );
  OAI22XL U5663 ( .A0(n4711), .A1(n360), .B0(n4720), .B1(n352), .Y(n1248) );
  OAI22XL U5664 ( .A0(n1145), .A1(n294), .B0(n1146), .B1(n286), .Y(n1138) );
  OAI22XL U5665 ( .A0(n4711), .A1(n358), .B0(n4720), .B1(n350), .Y(n1150) );
  OAI22XL U5666 ( .A0(n1145), .A1(n295), .B0(n1146), .B1(n287), .Y(n1203) );
  OAI22XL U5667 ( .A0(n4711), .A1(n359), .B0(n4720), .B1(n351), .Y(n1207) );
  OAI22XL U5668 ( .A0(n1167), .A1(n445), .B0(n1168), .B1(n437), .Y(n1473) );
  OAI22XL U5669 ( .A0(n1167), .A1(n444), .B0(n1168), .B1(n436), .Y(n1417) );
  OAI22XL U5670 ( .A0(n1167), .A1(n443), .B0(n1168), .B1(n435), .Y(n1376) );
  OAI22XL U5671 ( .A0(n1167), .A1(n442), .B0(n1168), .B1(n434), .Y(n1335) );
  OAI22XL U5672 ( .A0(n1167), .A1(n441), .B0(n1168), .B1(n433), .Y(n1294) );
  OAI22XL U5673 ( .A0(n1167), .A1(n440), .B0(n1168), .B1(n432), .Y(n1253) );
  OAI22XL U5674 ( .A0(n1167), .A1(n438), .B0(n1168), .B1(n430), .Y(n1163) );
  OAI22XL U5675 ( .A0(n1167), .A1(n439), .B0(n1168), .B1(n431), .Y(n1212) );
  OAI22XL U5676 ( .A0(n1080), .A1(n573), .B0(n4714), .B1(n565), .Y(n1426) );
  OAI22XL U5677 ( .A0(n1080), .A1(n572), .B0(n4714), .B1(n564), .Y(n1385) );
  OAI22XL U5678 ( .A0(n1080), .A1(n571), .B0(n4714), .B1(n563), .Y(n1344) );
  OAI22XL U5679 ( .A0(n1080), .A1(n570), .B0(n4714), .B1(n562), .Y(n1303) );
  OAI22XL U5680 ( .A0(n1080), .A1(n569), .B0(n4714), .B1(n561), .Y(n1262) );
  OAI22XL U5681 ( .A0(n1080), .A1(n568), .B0(n4714), .B1(n560), .Y(n1221) );
  OAI22XL U5682 ( .A0(n1080), .A1(n566), .B0(n4714), .B1(n558), .Y(n1076) );
  OAI22XL U5683 ( .A0(n1080), .A1(n567), .B0(n4714), .B1(n559), .Y(n1180) );
  OAI22XL U5684 ( .A0(n1169), .A1(n429), .B0(n4722), .B1(n421), .Y(n1472) );
  OAI22XL U5685 ( .A0(n1169), .A1(n428), .B0(n4722), .B1(n420), .Y(n1416) );
  OAI22XL U5686 ( .A0(n1169), .A1(n427), .B0(n4722), .B1(n419), .Y(n1375) );
  OAI22XL U5687 ( .A0(n1169), .A1(n426), .B0(n4722), .B1(n418), .Y(n1334) );
  OAI22XL U5688 ( .A0(n1169), .A1(n425), .B0(n4722), .B1(n417), .Y(n1293) );
  OAI22XL U5689 ( .A0(n1169), .A1(n424), .B0(n4722), .B1(n416), .Y(n1252) );
  OAI22XL U5690 ( .A0(n1169), .A1(n422), .B0(n4722), .B1(n414), .Y(n1162) );
  OAI22XL U5691 ( .A0(n1169), .A1(n423), .B0(n4722), .B1(n415), .Y(n1211) );
  OAI22XL U5692 ( .A0(n4707), .A1(n557), .B0(n1083), .B1(n549), .Y(n1425) );
  OAI22XL U5693 ( .A0(n4707), .A1(n556), .B0(n1083), .B1(n548), .Y(n1384) );
  OAI22XL U5694 ( .A0(n4707), .A1(n555), .B0(n1083), .B1(n547), .Y(n1343) );
  OAI22XL U5695 ( .A0(n4707), .A1(n554), .B0(n1083), .B1(n546), .Y(n1302) );
  OAI22XL U5696 ( .A0(n4707), .A1(n553), .B0(n1083), .B1(n545), .Y(n1261) );
  OAI22XL U5697 ( .A0(n4707), .A1(n552), .B0(n1083), .B1(n544), .Y(n1220) );
  OAI22XL U5698 ( .A0(n4707), .A1(n550), .B0(n1083), .B1(n542), .Y(n1075) );
  OAI22XL U5699 ( .A0(n4707), .A1(n551), .B0(n1083), .B1(n543), .Y(n1179) );
  OAI22XL U5700 ( .A0(n4716), .A1(n333), .B0(n1142), .B1(n325), .Y(n1464) );
  OAI22XL U5701 ( .A0(n1153), .A1(n397), .B0(n1154), .B1(n389), .Y(n1469) );
  OAI22XL U5702 ( .A0(n4716), .A1(n332), .B0(n1142), .B1(n324), .Y(n1410) );
  OAI22XL U5703 ( .A0(n1153), .A1(n396), .B0(n1154), .B1(n388), .Y(n1414) );
  OAI22XL U5704 ( .A0(n4716), .A1(n331), .B0(n1142), .B1(n323), .Y(n1369) );
  OAI22XL U5705 ( .A0(n1153), .A1(n395), .B0(n1154), .B1(n387), .Y(n1373) );
  OAI22XL U5706 ( .A0(n4716), .A1(n330), .B0(n1142), .B1(n322), .Y(n1328) );
  OAI22XL U5707 ( .A0(n1153), .A1(n394), .B0(n1154), .B1(n386), .Y(n1332) );
  OAI22XL U5708 ( .A0(n4716), .A1(n329), .B0(n1142), .B1(n321), .Y(n1287) );
  OAI22XL U5709 ( .A0(n1153), .A1(n393), .B0(n1154), .B1(n385), .Y(n1291) );
  OAI22XL U5710 ( .A0(n4716), .A1(n328), .B0(n1142), .B1(n320), .Y(n1246) );
  OAI22XL U5711 ( .A0(n1153), .A1(n392), .B0(n1154), .B1(n384), .Y(n1250) );
  OAI22XL U5712 ( .A0(n4716), .A1(n326), .B0(n1142), .B1(n318), .Y(n1140) );
  OAI22XL U5713 ( .A0(n1153), .A1(n390), .B0(n1154), .B1(n382), .Y(n1152) );
  OAI22XL U5714 ( .A0(n4716), .A1(n327), .B0(n1142), .B1(n319), .Y(n1205) );
  OAI22XL U5715 ( .A0(n1153), .A1(n391), .B0(n1154), .B1(n383), .Y(n1209) );
  OAI22XL U5716 ( .A0(n1165), .A1(n461), .B0(n1166), .B1(n453), .Y(n1474) );
  OAI22XL U5717 ( .A0(n1165), .A1(n460), .B0(n1166), .B1(n452), .Y(n1418) );
  OAI22XL U5718 ( .A0(n1165), .A1(n459), .B0(n1166), .B1(n451), .Y(n1377) );
  OAI22XL U5719 ( .A0(n1165), .A1(n458), .B0(n1166), .B1(n450), .Y(n1336) );
  OAI22XL U5720 ( .A0(n1165), .A1(n457), .B0(n1166), .B1(n449), .Y(n1295) );
  OAI22XL U5721 ( .A0(n1165), .A1(n456), .B0(n1166), .B1(n448), .Y(n1254) );
  OAI22XL U5722 ( .A0(n1165), .A1(n454), .B0(n1166), .B1(n446), .Y(n1164) );
  OAI22XL U5723 ( .A0(n1165), .A1(n455), .B0(n1166), .B1(n447), .Y(n1213) );
  OAI22XL U5724 ( .A0(n1078), .A1(n589), .B0(n1079), .B1(n581), .Y(n1427) );
  OAI22XL U5725 ( .A0(n1078), .A1(n588), .B0(n1079), .B1(n580), .Y(n1386) );
  OAI22XL U5726 ( .A0(n1078), .A1(n587), .B0(n1079), .B1(n579), .Y(n1345) );
  OAI22XL U5727 ( .A0(n1078), .A1(n586), .B0(n1079), .B1(n578), .Y(n1304) );
  OAI22XL U5728 ( .A0(n1078), .A1(n585), .B0(n1079), .B1(n577), .Y(n1263) );
  OAI22XL U5729 ( .A0(n1078), .A1(n584), .B0(n1079), .B1(n576), .Y(n1222) );
  OAI22XL U5730 ( .A0(n1078), .A1(n582), .B0(n1079), .B1(n574), .Y(n1077) );
  OAI22XL U5731 ( .A0(n1078), .A1(n583), .B0(n1079), .B1(n575), .Y(n1181) );
  AOI211XL U5732 ( .A0(n4069), .A1(n4749), .B0(n4076), .C0(reset), .Y(n4075)
         );
  OAI22XL U5733 ( .A0(n4685), .A1(n477), .B0(n1120), .B1(n469), .Y(n1447) );
  OAI22XL U5734 ( .A0(n4685), .A1(n476), .B0(n1120), .B1(n468), .Y(n1395) );
  OAI22XL U5735 ( .A0(n4685), .A1(n475), .B0(n1120), .B1(n467), .Y(n1354) );
  OAI22XL U5736 ( .A0(n4685), .A1(n474), .B0(n1120), .B1(n466), .Y(n1313) );
  OAI22XL U5737 ( .A0(n4685), .A1(n473), .B0(n1120), .B1(n465), .Y(n1272) );
  OAI22XL U5738 ( .A0(n4685), .A1(n472), .B0(n1120), .B1(n464), .Y(n1231) );
  OAI22XL U5739 ( .A0(n4685), .A1(n470), .B0(n1120), .B1(n462), .Y(n1109) );
  OAI22XL U5740 ( .A0(n4685), .A1(n471), .B0(n1120), .B1(n463), .Y(n1190) );
  OAI22XL U5741 ( .A0(n4687), .A1(n509), .B0(n4709), .B1(n501), .Y(n1449) );
  OAI22XL U5742 ( .A0(n4687), .A1(n508), .B0(n4709), .B1(n500), .Y(n1397) );
  OAI22XL U5743 ( .A0(n4687), .A1(n507), .B0(n4709), .B1(n499), .Y(n1356) );
  OAI22XL U5744 ( .A0(n4687), .A1(n506), .B0(n4709), .B1(n498), .Y(n1315) );
  OAI22XL U5745 ( .A0(n4687), .A1(n505), .B0(n4709), .B1(n497), .Y(n1274) );
  OAI22XL U5746 ( .A0(n4687), .A1(n504), .B0(n4709), .B1(n496), .Y(n1233) );
  OAI22XL U5747 ( .A0(n4687), .A1(n502), .B0(n4709), .B1(n494), .Y(n1111) );
  OAI22XL U5748 ( .A0(n4687), .A1(n503), .B0(n4709), .B1(n495), .Y(n1192) );
  OAI22XL U5749 ( .A0(n4715), .A1(n493), .B0(n4713), .B1(n485), .Y(n1448) );
  OAI22XL U5750 ( .A0(n4715), .A1(n492), .B0(n4713), .B1(n484), .Y(n1396) );
  OAI22XL U5751 ( .A0(n4715), .A1(n491), .B0(n4713), .B1(n483), .Y(n1355) );
  OAI22XL U5752 ( .A0(n4715), .A1(n490), .B0(n4713), .B1(n482), .Y(n1314) );
  OAI22XL U5753 ( .A0(n4715), .A1(n489), .B0(n4713), .B1(n481), .Y(n1273) );
  OAI22XL U5754 ( .A0(n4715), .A1(n488), .B0(n4713), .B1(n480), .Y(n1232) );
  OAI22XL U5755 ( .A0(n4715), .A1(n486), .B0(n4713), .B1(n478), .Y(n1110) );
  OAI22XL U5756 ( .A0(n4715), .A1(n487), .B0(n4713), .B1(n479), .Y(n1191) );
  OAI22XL U5757 ( .A0(n1113), .A1(n525), .B0(n1114), .B1(n517), .Y(n1450) );
  OAI22XL U5758 ( .A0(n1113), .A1(n524), .B0(n1114), .B1(n516), .Y(n1398) );
  OAI22XL U5759 ( .A0(n1113), .A1(n523), .B0(n1114), .B1(n515), .Y(n1357) );
  OAI22XL U5760 ( .A0(n1113), .A1(n522), .B0(n1114), .B1(n514), .Y(n1316) );
  OAI22XL U5761 ( .A0(n1113), .A1(n521), .B0(n1114), .B1(n513), .Y(n1275) );
  OAI22XL U5762 ( .A0(n1113), .A1(n520), .B0(n1114), .B1(n512), .Y(n1234) );
  OAI22XL U5763 ( .A0(n1113), .A1(n518), .B0(n1114), .B1(n510), .Y(n1112) );
  OAI22XL U5764 ( .A0(n1113), .A1(n519), .B0(n1114), .B1(n511), .Y(n1193) );
  CLKBUFX3 U5765 ( .A(cur_state), .Y(n5951) );
  NAND3X1 U5766 ( .A(n4060), .B(n963), .C(cmd_reg[2]), .Y(n4073) );
  CLKBUFX3 U5767 ( .A(cur_state), .Y(n5953) );
  CLKBUFX3 U5768 ( .A(cur_state), .Y(n5952) );
  CLKBUFX3 U5769 ( .A(n5785), .Y(n5784) );
  CLKBUFX3 U5770 ( .A(n5785), .Y(n5783) );
  CLKBUFX3 U5771 ( .A(n5785), .Y(n5782) );
  CLKBUFX3 U5772 ( .A(n5785), .Y(n5781) );
  CLKBUFX3 U5773 ( .A(n5444), .Y(n5452) );
  CLKBUFX3 U5774 ( .A(n5443), .Y(n5454) );
  CLKBUFX3 U5775 ( .A(n1052), .Y(n5787) );
  CLKBUFX3 U5776 ( .A(n1052), .Y(n5786) );
  CLKBUFX3 U5777 ( .A(n1052), .Y(n5790) );
  CLKBUFX3 U5778 ( .A(n5776), .Y(n5778) );
  CLKBUFX3 U5779 ( .A(n5450), .Y(n5444) );
  CLKBUFX3 U5780 ( .A(n5450), .Y(n5443) );
  CLKBUFX3 U5781 ( .A(n5851), .Y(n5854) );
  CLKBUFX3 U5782 ( .A(n5851), .Y(n5853) );
  CLKBUFX3 U5783 ( .A(n1022), .Y(n5852) );
  OAI22XL U5784 ( .A0(n5669), .A1(n5699), .B0(n3986), .B1(n5750), .Y(n4034) );
  OAI22XL U5785 ( .A0(n5669), .A1(n5695), .B0(n3986), .B1(n5746), .Y(n4026) );
  OAI22XL U5786 ( .A0(n5669), .A1(n5688), .B0(n3986), .B1(n5741), .Y(n4014) );
  OAI22XL U5787 ( .A0(n5669), .A1(n5684), .B0(n3986), .B1(n5737), .Y(n4008) );
  OAI22XL U5788 ( .A0(n5669), .A1(n5681), .B0(n3986), .B1(n5735), .Y(n4002) );
  OAI22XL U5789 ( .A0(n5669), .A1(n5675), .B0(n5728), .B1(n3986), .Y(n3984) );
  CLKBUFX3 U5790 ( .A(n1058), .Y(n5768) );
  CLKBUFX3 U5791 ( .A(n1058), .Y(n5769) );
  CLKBUFX3 U5792 ( .A(n1058), .Y(n5767) );
  CLKBUFX3 U5793 ( .A(n1058), .Y(n5770) );
  CLKBUFX3 U5794 ( .A(n1055), .Y(n5775) );
  CLKBUFX3 U5795 ( .A(n1058), .Y(n5771) );
  CLKBUFX3 U5796 ( .A(n5626), .Y(n5631) );
  CLKBUFX3 U5797 ( .A(n5246), .Y(n5249) );
  CLKBUFX3 U5798 ( .A(n5256), .Y(n5257) );
  CLKBUFX3 U5799 ( .A(n5256), .Y(n5258) );
  CLKBUFX3 U5800 ( .A(n5638), .Y(n5259) );
  CLKBUFX3 U5801 ( .A(n5626), .Y(n5630) );
  CLKBUFX3 U5802 ( .A(n5625), .Y(n5633) );
  CLKBUFX3 U5803 ( .A(n5266), .Y(n5642) );
  CLKBUFX3 U5804 ( .A(n5266), .Y(n5646) );
  CLKBUFX3 U5805 ( .A(n5256), .Y(n5643) );
  CLKBUFX3 U5806 ( .A(n5256), .Y(n5644) );
  CLKBUFX3 U5807 ( .A(n5256), .Y(n5645) );
  CLKBUFX3 U5808 ( .A(n5639), .Y(n5260) );
  CLKBUFX3 U5809 ( .A(n5639), .Y(n5261) );
  CLKBUFX3 U5810 ( .A(n5259), .Y(n5262) );
  CLKBUFX3 U5811 ( .A(n5640), .Y(n5264) );
  CLKBUFX3 U5812 ( .A(n5256), .Y(n5263) );
  CLKBUFX3 U5813 ( .A(n5624), .Y(n5635) );
  CLKBUFX3 U5814 ( .A(n5243), .Y(n5253) );
  CLKBUFX3 U5815 ( .A(n4749), .Y(n5265) );
  INVX4 U5816 ( .A(n5766), .Y(n5764) );
  INVX4 U5817 ( .A(n5766), .Y(n5765) );
  CLKBUFX3 U5818 ( .A(n1022), .Y(n5851) );
  NOR2BX2 U5819 ( .AN(n3980), .B(n4032), .Y(n3977) );
  OAI22XL U5820 ( .A0(n3980), .A1(n5695), .B0(n3981), .B1(n5746), .Y(n4025) );
  OAI22XL U5821 ( .A0(n3980), .A1(n5691), .B0(n3981), .B1(n5743), .Y(n4019) );
  OAI22XL U5822 ( .A0(n3980), .A1(n5688), .B0(n3981), .B1(n5740), .Y(n4013) );
  OAI22XL U5823 ( .A0(n3980), .A1(n5681), .B0(n3981), .B1(n5735), .Y(n4001) );
  OAI22XL U5824 ( .A0(n3980), .A1(n5675), .B0(n3981), .B1(n5728), .Y(n3979) );
  OAI22XL U5825 ( .A0(n3980), .A1(n5679), .B0(n3981), .B1(n5730), .Y(n3994) );
  OR3X2 U5826 ( .A(n6298), .B(n6270), .C(n6327), .Y(n4053) );
  CLKBUFX3 U5827 ( .A(n5442), .Y(n5433) );
  CLKBUFX3 U5828 ( .A(n5072), .Y(n5073) );
  CLKBUFX3 U5829 ( .A(n5637), .Y(n5627) );
  CLKBUFX3 U5830 ( .A(n5636), .Y(n5625) );
  CLKBUFX3 U5831 ( .A(n5076), .Y(n5438) );
  CLKBUFX3 U5832 ( .A(n5441), .Y(n5079) );
  CLKBUFX3 U5833 ( .A(n5636), .Y(n5624) );
  CLKBUFX3 U5834 ( .A(n5254), .Y(n5243) );
  INVX3 U5835 ( .A(n3370), .Y(n6512) );
  INVX3 U5836 ( .A(n3331), .Y(n6520) );
  INVX3 U5837 ( .A(n3292), .Y(n6528) );
  INVX3 U5838 ( .A(n3253), .Y(n6536) );
  INVX3 U5839 ( .A(n3214), .Y(n6544) );
  INVX3 U5840 ( .A(n3175), .Y(n6552) );
  INVX3 U5841 ( .A(n3136), .Y(n6560) );
  INVX3 U5842 ( .A(n3093), .Y(n6568) );
  INVX3 U5843 ( .A(n3053), .Y(n6513) );
  INVX3 U5844 ( .A(n3014), .Y(n6521) );
  INVX3 U5845 ( .A(n2975), .Y(n6529) );
  INVX3 U5846 ( .A(n2936), .Y(n6537) );
  INVX3 U5847 ( .A(n2897), .Y(n6545) );
  INVX3 U5848 ( .A(n2858), .Y(n6553) );
  INVX3 U5849 ( .A(n2819), .Y(n6561) );
  INVX3 U5850 ( .A(n2776), .Y(n6569) );
  INVX3 U5851 ( .A(n2102), .Y(n6516) );
  INVX3 U5852 ( .A(n2063), .Y(n6524) );
  INVX3 U5853 ( .A(n3648), .Y(n6519) );
  INVX3 U5854 ( .A(n3609), .Y(n6527) );
  INVX3 U5855 ( .A(n3570), .Y(n6535) );
  INVX3 U5856 ( .A(n2736), .Y(n6514) );
  INVX3 U5857 ( .A(n2697), .Y(n6522) );
  INVX3 U5858 ( .A(n2658), .Y(n6530) );
  INVX3 U5859 ( .A(n2619), .Y(n6538) );
  INVX3 U5860 ( .A(n2419), .Y(n6515) );
  INVX3 U5861 ( .A(n2380), .Y(n6523) );
  INVX3 U5862 ( .A(n2341), .Y(n6531) );
  INVX3 U5863 ( .A(n2302), .Y(n6539) );
  CLKINVX1 U5864 ( .A(n3727), .Y(n6566) );
  INVX3 U5865 ( .A(n3531), .Y(n6543) );
  INVX3 U5866 ( .A(n3492), .Y(n6551) );
  INVX3 U5867 ( .A(n3453), .Y(n6559) );
  INVX3 U5868 ( .A(n3410), .Y(n6567) );
  INVX3 U5869 ( .A(n2580), .Y(n6546) );
  INVX3 U5870 ( .A(n2541), .Y(n6554) );
  INVX3 U5871 ( .A(n2502), .Y(n6562) );
  INVX3 U5872 ( .A(n2459), .Y(n6570) );
  INVX3 U5873 ( .A(n2263), .Y(n6547) );
  INVX3 U5874 ( .A(n2224), .Y(n6555) );
  INVX3 U5875 ( .A(n2185), .Y(n6563) );
  INVX3 U5876 ( .A(n2142), .Y(n6571) );
  NOR3BXL U5877 ( .AN(n3358), .B(n6512), .C(n5818), .Y(n3361) );
  NOR3BXL U5878 ( .AN(n3319), .B(n6520), .C(n5817), .Y(n3322) );
  NOR3BXL U5879 ( .AN(n3280), .B(n6528), .C(n5817), .Y(n3283) );
  NOR3BXL U5880 ( .AN(n3241), .B(n6536), .C(n5817), .Y(n3244) );
  NOR3BXL U5881 ( .AN(n3202), .B(n6544), .C(n5817), .Y(n3205) );
  NOR3BXL U5882 ( .AN(n3163), .B(n6552), .C(n5817), .Y(n3166) );
  NOR3BXL U5883 ( .AN(n3124), .B(n6560), .C(n5817), .Y(n3127) );
  NOR3BXL U5884 ( .AN(n3080), .B(n6568), .C(n5817), .Y(n3083) );
  NOR3BXL U5885 ( .AN(n3041), .B(n6513), .C(n5817), .Y(n3044) );
  NOR3BXL U5886 ( .AN(n3002), .B(n6521), .C(n5817), .Y(n3005) );
  NOR3BXL U5887 ( .AN(n2963), .B(n6529), .C(n5817), .Y(n2966) );
  NOR3BXL U5888 ( .AN(n2924), .B(n6537), .C(n5816), .Y(n2927) );
  NOR3BXL U5889 ( .AN(n2885), .B(n6545), .C(n5816), .Y(n2888) );
  NOR3BXL U5890 ( .AN(n2846), .B(n6553), .C(n5816), .Y(n2849) );
  NOR3BXL U5891 ( .AN(n2807), .B(n6561), .C(n5816), .Y(n2810) );
  NOR3BXL U5892 ( .AN(n2763), .B(n6569), .C(n5816), .Y(n2766) );
  NOR3BXL U5893 ( .AN(n2090), .B(n6516), .C(n5817), .Y(n2093) );
  NOR3BXL U5894 ( .AN(n2051), .B(n6524), .C(n5815), .Y(n2054) );
  NOR3BXL U5895 ( .AN(n4041), .B(n6510), .C(n5817), .Y(n4044) );
  NOR3BXL U5896 ( .AN(n3953), .B(n6518), .C(n5819), .Y(n3956) );
  NOR3BXL U5897 ( .AN(n3914), .B(n6526), .C(n5819), .Y(n3917) );
  NOR3BXL U5898 ( .AN(n3875), .B(n6534), .C(n5818), .Y(n3878) );
  NOR3BXL U5899 ( .AN(n3675), .B(n6511), .C(n5818), .Y(n3678) );
  NOR3BXL U5900 ( .AN(n3636), .B(n6519), .C(n5818), .Y(n3639) );
  NOR3BXL U5901 ( .AN(n3597), .B(n6527), .C(n5818), .Y(n3600) );
  NOR3BXL U5902 ( .AN(n3558), .B(n6535), .C(n5818), .Y(n3561) );
  NOR3BXL U5903 ( .AN(n2724), .B(n6514), .C(n5816), .Y(n2727) );
  NOR3BXL U5904 ( .AN(n2685), .B(n6522), .C(n5816), .Y(n2688) );
  NOR3BXL U5905 ( .AN(n2646), .B(n6530), .C(n5816), .Y(n2649) );
  NOR3BXL U5906 ( .AN(n2607), .B(n6538), .C(n5816), .Y(n2610) );
  NOR3BXL U5907 ( .AN(n2407), .B(n6515), .C(n5817), .Y(n2410) );
  NOR3BXL U5908 ( .AN(n2368), .B(n6523), .C(n5817), .Y(n2371) );
  NOR3BXL U5909 ( .AN(n2329), .B(n6531), .C(n5817), .Y(n2332) );
  NOR3BXL U5910 ( .AN(n2290), .B(n6539), .C(n5817), .Y(n2293) );
  NOR3BXL U5911 ( .AN(n3836), .B(n6542), .C(n5818), .Y(n3839) );
  NOR3BXL U5912 ( .AN(n3797), .B(n6550), .C(n5819), .Y(n3800) );
  NOR3BXL U5913 ( .AN(n3758), .B(n6558), .C(n5818), .Y(n3761) );
  NOR3BXL U5914 ( .AN(n3714), .B(n6566), .C(n5818), .Y(n3717) );
  NOR3BXL U5915 ( .AN(n3519), .B(n6543), .C(n5818), .Y(n3522) );
  NOR3BXL U5916 ( .AN(n3480), .B(n6551), .C(n5818), .Y(n3483) );
  NOR3BXL U5917 ( .AN(n3441), .B(n6559), .C(n5818), .Y(n3444) );
  NOR3BXL U5918 ( .AN(n3397), .B(n6567), .C(n5817), .Y(n3400) );
  NOR3BXL U5919 ( .AN(n2568), .B(n6546), .C(n5816), .Y(n2571) );
  NOR3BXL U5920 ( .AN(n2529), .B(n6554), .C(n5816), .Y(n2532) );
  NOR3BXL U5921 ( .AN(n2490), .B(n6562), .C(n5816), .Y(n2493) );
  NOR3BXL U5922 ( .AN(n2446), .B(n6570), .C(n5817), .Y(n2449) );
  NOR3BXL U5923 ( .AN(n2251), .B(n6547), .C(n5817), .Y(n2254) );
  NOR3BXL U5924 ( .AN(n2212), .B(n6555), .C(n5817), .Y(n2215) );
  NOR3BXL U5925 ( .AN(n2173), .B(n6563), .C(n5816), .Y(n2176) );
  NOR3BXL U5926 ( .AN(n2129), .B(n6571), .C(n5818), .Y(n2132) );
  CLKBUFX3 U5927 ( .A(n5076), .Y(n5440) );
  CLKBUFX3 U5928 ( .A(n5070), .Y(n5081) );
  CLKBUFX3 U5929 ( .A(n5727), .Y(n5728) );
  CLKBUFX3 U5930 ( .A(n5749), .Y(n5750) );
  CLKBUFX3 U5931 ( .A(n5734), .Y(n5735) );
  INVX3 U5932 ( .A(n1027), .Y(n6573) );
  INVX3 U5933 ( .A(n1771), .Y(n6517) );
  INVX3 U5934 ( .A(n1727), .Y(n6525) );
  INVX3 U5935 ( .A(n1683), .Y(n6533) );
  INVX3 U5936 ( .A(n1639), .Y(n6541) );
  INVX3 U5937 ( .A(n1595), .Y(n6549) );
  INVX3 U5938 ( .A(n1551), .Y(n6557) );
  INVX3 U5939 ( .A(n1507), .Y(n6565) );
  INVX3 U5940 ( .A(n2016), .Y(n6532) );
  INVX3 U5941 ( .A(n1977), .Y(n6540) );
  INVX3 U5942 ( .A(n1938), .Y(n6548) );
  INVX3 U5943 ( .A(n1899), .Y(n6556) );
  INVX3 U5944 ( .A(n1860), .Y(n6564) );
  INVX3 U5945 ( .A(n1816), .Y(n6572) );
  NOR3BXL U5946 ( .AN(n1033), .B(n6573), .C(n5817), .Y(n1026) );
  CLKBUFX3 U5947 ( .A(n5698), .Y(n5699) );
  CLKBUFX3 U5948 ( .A(n6422), .Y(n5695) );
  CLKBUFX3 U5949 ( .A(n6421), .Y(n5691) );
  CLKBUFX3 U5950 ( .A(n6420), .Y(n5688) );
  CLKBUFX3 U5951 ( .A(n6419), .Y(n5684) );
  CLKBUFX3 U5952 ( .A(n5750), .Y(n5751) );
  CLKBUFX3 U5953 ( .A(n5747), .Y(n5748) );
  CLKBUFX3 U5954 ( .A(n5746), .Y(n5747) );
  CLKBUFX3 U5955 ( .A(n6507), .Y(n5744) );
  CLKBUFX3 U5956 ( .A(n5744), .Y(n5745) );
  CLKBUFX3 U5957 ( .A(n6257), .Y(n5741) );
  CLKBUFX3 U5958 ( .A(n5738), .Y(n5739) );
  CLKBUFX3 U5959 ( .A(n5737), .Y(n5738) );
  CLKBUFX3 U5960 ( .A(n5733), .Y(n5736) );
  CLKBUFX3 U5961 ( .A(n5728), .Y(n5729) );
  CLKBUFX3 U5962 ( .A(n5730), .Y(n5732) );
  AND3X2 U5963 ( .A(n2010), .B(n2016), .C(n5824), .Y(n2012) );
  AND3X2 U5964 ( .A(n1971), .B(n1977), .C(n5824), .Y(n1973) );
  AND3X2 U5965 ( .A(n1932), .B(n1938), .C(n5826), .Y(n1934) );
  AND3X2 U5966 ( .A(n1810), .B(n1816), .C(n5825), .Y(n1812) );
  CLKBUFX3 U5967 ( .A(n6007), .Y(n5675) );
  CLKBUFX3 U5968 ( .A(n5678), .Y(n5679) );
  CLKBUFX3 U5969 ( .A(n5698), .Y(n5700) );
  CLKBUFX3 U5970 ( .A(n5700), .Y(n5701) );
  CLKBUFX3 U5971 ( .A(n5696), .Y(n5697) );
  CLKBUFX3 U5972 ( .A(n6003), .Y(n5696) );
  CLKBUFX3 U5973 ( .A(n5692), .Y(n5694) );
  CLKBUFX3 U5974 ( .A(n6421), .Y(n5692) );
  CLKBUFX3 U5975 ( .A(n5692), .Y(n5693) );
  CLKBUFX3 U5976 ( .A(n5688), .Y(n5689) );
  CLKBUFX3 U5977 ( .A(n5689), .Y(n5690) );
  CLKBUFX3 U5978 ( .A(n5685), .Y(n5687) );
  CLKBUFX3 U5979 ( .A(n6419), .Y(n5685) );
  CLKBUFX3 U5980 ( .A(n5685), .Y(n5686) );
  CLKBUFX3 U5981 ( .A(n5682), .Y(n5683) );
  CLKBUFX3 U5982 ( .A(n5681), .Y(n5682) );
  CLKBUFX3 U5983 ( .A(n5676), .Y(n5677) );
  CLKBUFX3 U5984 ( .A(n6070), .Y(n5676) );
  CLKBUFX3 U5985 ( .A(n5679), .Y(n5680) );
  CLKBUFX3 U5986 ( .A(n4827), .Y(n5766) );
  NOR2X1 U5987 ( .A(n5845), .B(n5831), .Y(n1022) );
  CLKBUFX3 U5988 ( .A(n6502), .Y(n5724) );
  CLKBUFX3 U5989 ( .A(n6502), .Y(n5725) );
  CLKBUFX3 U5990 ( .A(n6502), .Y(n5726) );
  CLKBUFX3 U5991 ( .A(n6131), .Y(n5721) );
  CLKBUFX3 U5992 ( .A(n4817), .Y(n5722) );
  CLKBUFX3 U5993 ( .A(n6098), .Y(n5723) );
  CLKBUFX3 U5994 ( .A(n6501), .Y(n5718) );
  CLKBUFX3 U5995 ( .A(n6501), .Y(n5719) );
  CLKBUFX3 U5996 ( .A(n6501), .Y(n5720) );
  CLKBUFX3 U5997 ( .A(n6162), .Y(n5715) );
  CLKBUFX3 U5998 ( .A(n6132), .Y(n5716) );
  CLKBUFX3 U5999 ( .A(n6132), .Y(n5717) );
  CLKBUFX3 U6000 ( .A(n5711), .Y(n5712) );
  CLKBUFX3 U6001 ( .A(n5711), .Y(n5713) );
  CLKBUFX3 U6002 ( .A(n5711), .Y(n5714) );
  CLKBUFX3 U6003 ( .A(n6500), .Y(n5708) );
  CLKBUFX3 U6004 ( .A(n6500), .Y(n5709) );
  CLKBUFX3 U6005 ( .A(n6500), .Y(n5710) );
  CLKBUFX3 U6006 ( .A(n6165), .Y(n5702) );
  CLKBUFX3 U6007 ( .A(n6165), .Y(n5703) );
  CLKBUFX3 U6008 ( .A(n6101), .Y(n5704) );
  CLKBUFX3 U6009 ( .A(n6133), .Y(n5705) );
  CLKBUFX3 U6010 ( .A(n6100), .Y(n5706) );
  CLKBUFX3 U6011 ( .A(n6100), .Y(n5707) );
  CLKINVX1 U6012 ( .A(n6204), .Y(n6229) );
  OA22X2 U6013 ( .A0(n2014), .A1(n5772), .B0(n5770), .B1(n2010), .Y(n2025) );
  OAI221XL U6014 ( .A0(n5777), .A1(n4040), .B0(n4664), .B1(n4054), .C0(n4055), 
        .Y(n4049) );
  OAI221XL U6015 ( .A0(n5780), .A1(n3713), .B0(n4660), .B1(n3727), .C0(n3728), 
        .Y(n3723) );
  OAI221X1 U6016 ( .A0(n5780), .A1(n3518), .B0(n4658), .B1(n3531), .C0(n3532), 
        .Y(n3527) );
  OAI221X1 U6017 ( .A0(n5780), .A1(n3479), .B0(n4659), .B1(n3492), .C0(n3493), 
        .Y(n3488) );
  OAI221X1 U6018 ( .A0(n5780), .A1(n3440), .B0(n4663), .B1(n3453), .C0(n3454), 
        .Y(n3449) );
  OAI221X1 U6019 ( .A0(n5780), .A1(n3396), .B0(n4661), .B1(n3410), .C0(n3411), 
        .Y(n3406) );
  OAI221X1 U6020 ( .A0(n5780), .A1(n3357), .B0(n4664), .B1(n3370), .C0(n3371), 
        .Y(n3366) );
  OAI221X1 U6021 ( .A0(n5780), .A1(n3318), .B0(n4663), .B1(n3331), .C0(n3332), 
        .Y(n3327) );
  OAI221X1 U6022 ( .A0(n5780), .A1(n3279), .B0(n4657), .B1(n3292), .C0(n3293), 
        .Y(n3288) );
  OA22X2 U6023 ( .A0(n3247), .A1(n5773), .B0(n5767), .B1(n3241), .Y(n3254) );
  OAI221X1 U6024 ( .A0(n5779), .A1(n3201), .B0(n4665), .B1(n3214), .C0(n3215), 
        .Y(n3210) );
  OAI221X1 U6025 ( .A0(n5779), .A1(n3162), .B0(n4659), .B1(n3175), .C0(n3176), 
        .Y(n3171) );
  OA22X2 U6026 ( .A0(n3169), .A1(n5772), .B0(n5767), .B1(n3163), .Y(n3176) );
  OA22X2 U6027 ( .A0(n3130), .A1(n5773), .B0(n5767), .B1(n3124), .Y(n3137) );
  OA22X2 U6028 ( .A0(n3086), .A1(n5773), .B0(n5767), .B1(n3080), .Y(n3094) );
  OAI221X1 U6029 ( .A0(n5779), .A1(n3040), .B0(n4657), .B1(n3053), .C0(n3054), 
        .Y(n3049) );
  OAI221X1 U6030 ( .A0(n5779), .A1(n3001), .B0(n4657), .B1(n3014), .C0(n3015), 
        .Y(n3010) );
  OAI221X1 U6031 ( .A0(n5779), .A1(n2962), .B0(n4657), .B1(n2975), .C0(n2976), 
        .Y(n2971) );
  OAI221X1 U6032 ( .A0(n5779), .A1(n2923), .B0(n4664), .B1(n2936), .C0(n2937), 
        .Y(n2932) );
  OAI221X1 U6033 ( .A0(n5779), .A1(n2884), .B0(n4659), .B1(n2897), .C0(n2898), 
        .Y(n2893) );
  OA22X2 U6034 ( .A0(n2891), .A1(n5773), .B0(n5768), .B1(n2885), .Y(n2898) );
  OAI221X1 U6035 ( .A0(n5779), .A1(n2845), .B0(n4658), .B1(n2858), .C0(n2859), 
        .Y(n2854) );
  OA22X2 U6036 ( .A0(n2852), .A1(n5773), .B0(n5768), .B1(n2846), .Y(n2859) );
  OAI221X1 U6037 ( .A0(n5779), .A1(n2806), .B0(n4665), .B1(n2819), .C0(n2820), 
        .Y(n2815) );
  OAI221X1 U6038 ( .A0(n5779), .A1(n2762), .B0(n4665), .B1(n2776), .C0(n2777), 
        .Y(n2772) );
  OAI221X1 U6039 ( .A0(n5779), .A1(n2684), .B0(n4657), .B1(n2697), .C0(n2698), 
        .Y(n2693) );
  OA22X2 U6040 ( .A0(n2691), .A1(n5773), .B0(n5768), .B1(n2685), .Y(n2698) );
  OAI221X1 U6041 ( .A0(n5778), .A1(n2645), .B0(n4658), .B1(n2658), .C0(n2659), 
        .Y(n2654) );
  OAI221X1 U6042 ( .A0(n5778), .A1(n2606), .B0(n4659), .B1(n2619), .C0(n2620), 
        .Y(n2615) );
  OA22X2 U6043 ( .A0(n2613), .A1(n5773), .B0(n5768), .B1(n2607), .Y(n2620) );
  OAI221X1 U6044 ( .A0(n5778), .A1(n2406), .B0(n4659), .B1(n2419), .C0(n2420), 
        .Y(n2415) );
  OAI221X1 U6045 ( .A0(n5778), .A1(n2367), .B0(n4661), .B1(n2380), .C0(n2381), 
        .Y(n2376) );
  OAI221X1 U6046 ( .A0(n5778), .A1(n2328), .B0(n4661), .B1(n2341), .C0(n2342), 
        .Y(n2337) );
  OAI221X1 U6047 ( .A0(n5778), .A1(n2289), .B0(n4663), .B1(n2302), .C0(n2303), 
        .Y(n2298) );
  OA22X2 U6048 ( .A0(n2296), .A1(n5773), .B0(n5769), .B1(n2290), .Y(n2303) );
  OAI221X1 U6049 ( .A0(n5778), .A1(n2089), .B0(n4663), .B1(n2102), .C0(n2103), 
        .Y(n2098) );
  OAI221X1 U6050 ( .A0(n5778), .A1(n2567), .B0(n4665), .B1(n2580), .C0(n2581), 
        .Y(n2576) );
  OAI221X1 U6051 ( .A0(n5778), .A1(n2528), .B0(n4665), .B1(n2541), .C0(n2542), 
        .Y(n2537) );
  OAI221X1 U6052 ( .A0(n5778), .A1(n2489), .B0(n4663), .B1(n2502), .C0(n2503), 
        .Y(n2498) );
  OAI221X1 U6053 ( .A0(n5778), .A1(n2445), .B0(n4665), .B1(n2459), .C0(n2460), 
        .Y(n2455) );
  OA22X2 U6054 ( .A0(n2452), .A1(n5773), .B0(n5769), .B1(n2446), .Y(n2460) );
  OAI221X1 U6055 ( .A0(n5778), .A1(n2250), .B0(n4664), .B1(n2263), .C0(n2264), 
        .Y(n2259) );
  OA22X2 U6056 ( .A0(n2257), .A1(n5773), .B0(n5769), .B1(n2251), .Y(n2264) );
  OAI221X1 U6057 ( .A0(n5778), .A1(n2211), .B0(n4657), .B1(n2224), .C0(n2225), 
        .Y(n2220) );
  OAI221X1 U6058 ( .A0(n5778), .A1(n2172), .B0(n4660), .B1(n2185), .C0(n2186), 
        .Y(n2181) );
  OAI221X1 U6059 ( .A0(n5778), .A1(n2128), .B0(n4664), .B1(n2142), .C0(n2143), 
        .Y(n2138) );
  AOI221XL U6060 ( .A0(n6631), .A1(n4696), .B0(n6566), .B1(n4649), .C0(n3726), 
        .Y(n3725) );
  OAI22XL U6061 ( .A0(n5786), .A1(n3714), .B0(n5783), .B1(n3720), .Y(n3726) );
  AOI221X1 U6062 ( .A0(n6616), .A1(n4696), .B0(n6551), .B1(n4650), .C0(n3491), 
        .Y(n3490) );
  OAI22X2 U6063 ( .A0(n5787), .A1(n3480), .B0(n5785), .B1(n3486), .Y(n3491) );
  AOI221X1 U6064 ( .A0(n6624), .A1(n4696), .B0(n6559), .B1(n4650), .C0(n3452), 
        .Y(n3451) );
  OAI22X2 U6065 ( .A0(n5787), .A1(n3441), .B0(n5785), .B1(n3447), .Y(n3452) );
  AOI221X1 U6066 ( .A0(n6632), .A1(n4696), .B0(n6567), .B1(n4650), .C0(n3409), 
        .Y(n3408) );
  OAI22X2 U6067 ( .A0(n5787), .A1(n3397), .B0(n5785), .B1(n3403), .Y(n3409) );
  AOI221X1 U6068 ( .A0(n6577), .A1(n4696), .B0(n6512), .B1(n4650), .C0(n3369), 
        .Y(n3368) );
  OAI22X2 U6069 ( .A0(n5787), .A1(n3358), .B0(n5785), .B1(n3364), .Y(n3369) );
  AOI221X1 U6070 ( .A0(n6585), .A1(n4696), .B0(n6520), .B1(n4650), .C0(n3330), 
        .Y(n3329) );
  OAI22X2 U6071 ( .A0(n5787), .A1(n3319), .B0(n5785), .B1(n3325), .Y(n3330) );
  AOI221X1 U6072 ( .A0(n6593), .A1(n4696), .B0(n6528), .B1(n4650), .C0(n3291), 
        .Y(n3290) );
  OAI22X2 U6073 ( .A0(n5787), .A1(n3280), .B0(n5785), .B1(n3286), .Y(n3291) );
  AOI221X1 U6074 ( .A0(n6601), .A1(n4696), .B0(n6536), .B1(n4650), .C0(n3252), 
        .Y(n3251) );
  OAI22X2 U6075 ( .A0(n5787), .A1(n3241), .B0(n5785), .B1(n3247), .Y(n3252) );
  AOI221X1 U6076 ( .A0(n6609), .A1(n4696), .B0(n6544), .B1(n4650), .C0(n3213), 
        .Y(n3212) );
  OAI22X2 U6077 ( .A0(n5787), .A1(n3202), .B0(n5785), .B1(n3208), .Y(n3213) );
  OAI22X1 U6078 ( .A0(n5787), .A1(n3163), .B0(n5785), .B1(n3169), .Y(n3174) );
  OAI22X1 U6079 ( .A0(n5787), .A1(n3124), .B0(n5785), .B1(n3130), .Y(n3135) );
  OAI22X1 U6080 ( .A0(n5787), .A1(n3080), .B0(n5785), .B1(n3086), .Y(n3092) );
  OAI22X1 U6081 ( .A0(n5787), .A1(n3041), .B0(n5785), .B1(n3047), .Y(n3052) );
  OAI22X1 U6082 ( .A0(n5787), .A1(n3002), .B0(n5785), .B1(n3008), .Y(n3013) );
  AOI221X1 U6083 ( .A0(n6594), .A1(n4696), .B0(n6529), .B1(n4650), .C0(n2974), 
        .Y(n2973) );
  AOI221X1 U6084 ( .A0(n6602), .A1(n4696), .B0(n6537), .B1(n4650), .C0(n2935), 
        .Y(n2934) );
  OAI22X2 U6085 ( .A0(n4645), .A1(n2924), .B0(n5785), .B1(n2930), .Y(n2935) );
  AOI221X1 U6086 ( .A0(n6610), .A1(n4696), .B0(n6545), .B1(n4650), .C0(n2896), 
        .Y(n2895) );
  OAI22X2 U6087 ( .A0(n4645), .A1(n2885), .B0(n5785), .B1(n2891), .Y(n2896) );
  AOI221X1 U6088 ( .A0(n6618), .A1(n4696), .B0(n6553), .B1(n4650), .C0(n2857), 
        .Y(n2856) );
  OAI22X2 U6089 ( .A0(n4645), .A1(n2846), .B0(n5785), .B1(n2852), .Y(n2857) );
  AOI221X1 U6090 ( .A0(n6626), .A1(n4696), .B0(n6561), .B1(n4650), .C0(n2818), 
        .Y(n2817) );
  OAI22X2 U6091 ( .A0(n4645), .A1(n2807), .B0(n5785), .B1(n2813), .Y(n2818) );
  AOI221X1 U6092 ( .A0(n6634), .A1(n4696), .B0(n6569), .B1(n4650), .C0(n2775), 
        .Y(n2774) );
  OAI22X2 U6093 ( .A0(n4645), .A1(n2763), .B0(n5785), .B1(n2769), .Y(n2775) );
  AOI221X1 U6094 ( .A0(n6579), .A1(n4696), .B0(n6514), .B1(n4650), .C0(n2735), 
        .Y(n2734) );
  OAI22X2 U6095 ( .A0(n4645), .A1(n2724), .B0(n5785), .B1(n2730), .Y(n2735) );
  AOI221X1 U6096 ( .A0(n6587), .A1(n4696), .B0(n6522), .B1(n4649), .C0(n2696), 
        .Y(n2695) );
  OAI22X2 U6097 ( .A0(n4645), .A1(n2685), .B0(n5785), .B1(n2691), .Y(n2696) );
  OAI22X1 U6098 ( .A0(n4645), .A1(n2646), .B0(n5785), .B1(n2652), .Y(n2657) );
  OAI22X1 U6099 ( .A0(n4645), .A1(n2607), .B0(n5785), .B1(n2613), .Y(n2618) );
  OAI22X1 U6100 ( .A0(n4645), .A1(n2568), .B0(n5785), .B1(n2574), .Y(n2579) );
  OAI22X1 U6101 ( .A0(n4645), .A1(n2529), .B0(n5785), .B1(n2535), .Y(n2540) );
  OAI22X1 U6102 ( .A0(n4645), .A1(n2490), .B0(n5785), .B1(n2496), .Y(n2501) );
  AOI221X1 U6103 ( .A0(n6635), .A1(n4696), .B0(n6570), .B1(n4649), .C0(n2458), 
        .Y(n2457) );
  AOI221X1 U6104 ( .A0(n6580), .A1(n4696), .B0(n6515), .B1(n4650), .C0(n2418), 
        .Y(n2417) );
  AOI221X1 U6105 ( .A0(n6588), .A1(n4696), .B0(n6523), .B1(n4650), .C0(n2379), 
        .Y(n2378) );
  AOI221X1 U6106 ( .A0(n6596), .A1(n4696), .B0(n6531), .B1(n4650), .C0(n2340), 
        .Y(n2339) );
  AOI221X1 U6107 ( .A0(n6604), .A1(n4696), .B0(n6539), .B1(n4649), .C0(n2301), 
        .Y(n2300) );
  AOI221X1 U6108 ( .A0(n6612), .A1(n4696), .B0(n6547), .B1(n4649), .C0(n2262), 
        .Y(n2261) );
  AOI221X1 U6109 ( .A0(n6620), .A1(n4696), .B0(n6555), .B1(n4650), .C0(n2223), 
        .Y(n2222) );
  AOI221X1 U6110 ( .A0(n6628), .A1(n4696), .B0(n6563), .B1(n4650), .C0(n2184), 
        .Y(n2183) );
  OAI22X1 U6111 ( .A0(n4638), .A1(n2010), .B0(n5785), .B1(n2014), .Y(n2024) );
  AOI211X1 U6112 ( .A0(n6323), .A1(n6334), .B0(n6322), .C0(n6337), .Y(n6324)
         );
  AOI31X1 U6113 ( .A0(n6259), .A1(n6238), .A2(n6253), .B0(n6256), .Y(n6239) );
  OAI22X1 U6114 ( .A0(n5913), .A1(n1033), .B0(n1047), .B1(n4637), .Y(n1046) );
  AOI221X1 U6115 ( .A0(n6638), .A1(n4696), .B0(n6573), .B1(n4649), .C0(n1051), 
        .Y(n1047) );
  OAI22X2 U6116 ( .A0(n5790), .A1(n1033), .B0(n1032), .B1(n5785), .Y(n1051) );
  CLKINVX1 U6117 ( .A(n4829), .Y(n4894) );
  CLKBUFX3 U6118 ( .A(n5955), .Y(n5650) );
  CLKBUFX3 U6119 ( .A(n5955), .Y(n5649) );
  CLKBUFX3 U6120 ( .A(n5956), .Y(n5272) );
  CLKBUFX3 U6121 ( .A(n4893), .Y(n5271) );
  CLKINVX1 U6122 ( .A(n5955), .Y(n4893) );
  CLKBUFX3 U6123 ( .A(n5071), .Y(n5070) );
  AOI222X4 U6124 ( .A0(n5831), .A1(n4042), .B0(n4040), .B1(n4043), .C0(n5846), 
        .C1(n6510), .Y(n3988) );
  AO21X1 U6125 ( .A0(n5799), .A1(n6510), .B0(n4044), .Y(n4043) );
  AOI222X4 U6126 ( .A0(n5831), .A1(n3954), .B0(n3952), .B1(n3955), .C0(n5848), 
        .C1(n6518), .Y(n3934) );
  AO21X1 U6127 ( .A0(n5802), .A1(n6518), .B0(n3956), .Y(n3955) );
  AOI222X4 U6128 ( .A0(n5831), .A1(n3915), .B0(n3913), .B1(n3916), .C0(n5848), 
        .C1(n6526), .Y(n3895) );
  AO21X1 U6129 ( .A0(n5801), .A1(n6526), .B0(n3917), .Y(n3916) );
  AOI222X4 U6130 ( .A0(n5831), .A1(n3876), .B0(n3874), .B1(n3877), .C0(n5848), 
        .C1(n6534), .Y(n3856) );
  AO21X1 U6131 ( .A0(n5803), .A1(n6534), .B0(n3878), .Y(n3877) );
  AOI222X4 U6132 ( .A0(n5831), .A1(n3676), .B0(n3674), .B1(n3677), .C0(n5848), 
        .C1(n6511), .Y(n3656) );
  AO21X1 U6133 ( .A0(n5803), .A1(n6511), .B0(n3678), .Y(n3677) );
  AOI222X4 U6134 ( .A0(n5831), .A1(n3637), .B0(n3635), .B1(n3638), .C0(n5848), 
        .C1(n6519), .Y(n3617) );
  AO21X1 U6135 ( .A0(n5801), .A1(n6519), .B0(n3639), .Y(n3638) );
  AOI222X4 U6136 ( .A0(n5832), .A1(n3598), .B0(n3596), .B1(n3599), .C0(n5848), 
        .C1(n6527), .Y(n3578) );
  AO21X1 U6137 ( .A0(n5806), .A1(n6527), .B0(n3600), .Y(n3599) );
  AOI222X4 U6138 ( .A0(n5832), .A1(n3559), .B0(n3557), .B1(n3560), .C0(n5848), 
        .C1(n6535), .Y(n3539) );
  AO21X1 U6139 ( .A0(n5806), .A1(n6535), .B0(n3561), .Y(n3560) );
  AOI222X4 U6140 ( .A0(n5833), .A1(n2725), .B0(n2723), .B1(n2726), .C0(n5847), 
        .C1(n6514), .Y(n2705) );
  AO21X1 U6141 ( .A0(n5805), .A1(n6514), .B0(n2727), .Y(n2726) );
  AOI222X4 U6142 ( .A0(n5831), .A1(n2686), .B0(n2684), .B1(n2687), .C0(n5846), 
        .C1(n6522), .Y(n2666) );
  AO21X1 U6143 ( .A0(n5805), .A1(n6522), .B0(n2688), .Y(n2687) );
  AOI222X4 U6144 ( .A0(n5832), .A1(n2647), .B0(n2645), .B1(n2648), .C0(n5846), 
        .C1(n6530), .Y(n2627) );
  AO21X1 U6145 ( .A0(n5805), .A1(n6530), .B0(n2649), .Y(n2648) );
  AOI222X4 U6146 ( .A0(n5832), .A1(n2608), .B0(n2606), .B1(n2609), .C0(n5846), 
        .C1(n6538), .Y(n2588) );
  AO21X1 U6147 ( .A0(n5805), .A1(n6538), .B0(n2610), .Y(n2609) );
  AOI222X4 U6148 ( .A0(n5832), .A1(n2408), .B0(n2406), .B1(n2409), .C0(n5846), 
        .C1(n6515), .Y(n2388) );
  AO21X1 U6149 ( .A0(n5805), .A1(n6515), .B0(n2410), .Y(n2409) );
  AOI222X4 U6150 ( .A0(n5832), .A1(n2369), .B0(n2367), .B1(n2370), .C0(n5846), 
        .C1(n6523), .Y(n2349) );
  AO21X1 U6151 ( .A0(n5805), .A1(n6523), .B0(n2371), .Y(n2370) );
  AOI222X4 U6152 ( .A0(n5832), .A1(n2330), .B0(n2328), .B1(n2331), .C0(n5846), 
        .C1(n6531), .Y(n2310) );
  AO21X1 U6153 ( .A0(n5805), .A1(n6531), .B0(n2332), .Y(n2331) );
  AOI222X4 U6154 ( .A0(n5831), .A1(n2291), .B0(n2289), .B1(n2292), .C0(n5846), 
        .C1(n6539), .Y(n2271) );
  AO21X1 U6155 ( .A0(n5805), .A1(n6539), .B0(n2293), .Y(n2292) );
  NAND2X1 U6156 ( .A(n3096), .B(n1783), .Y(n3370) );
  NAND2X1 U6157 ( .A(n3096), .B(n1738), .Y(n3331) );
  NAND2X1 U6158 ( .A(n3096), .B(n1694), .Y(n3292) );
  NAND2X1 U6159 ( .A(n3096), .B(n1650), .Y(n3253) );
  NAND2X1 U6160 ( .A(n3096), .B(n1606), .Y(n3214) );
  NAND2X1 U6161 ( .A(n3096), .B(n1562), .Y(n3175) );
  NAND2X1 U6162 ( .A(n3096), .B(n1518), .Y(n3136) );
  NAND2X1 U6163 ( .A(n3096), .B(n1062), .Y(n3093) );
  NAND2X1 U6164 ( .A(n2779), .B(n1783), .Y(n3053) );
  NAND2X1 U6165 ( .A(n2779), .B(n1738), .Y(n3014) );
  NAND2X1 U6166 ( .A(n2779), .B(n1694), .Y(n2975) );
  NAND2X1 U6167 ( .A(n2779), .B(n1650), .Y(n2936) );
  NAND2X1 U6168 ( .A(n2779), .B(n1606), .Y(n2897) );
  NAND2X1 U6169 ( .A(n2779), .B(n1562), .Y(n2858) );
  NAND2X1 U6170 ( .A(n2779), .B(n1518), .Y(n2819) );
  NAND2X1 U6171 ( .A(n2779), .B(n1062), .Y(n2776) );
  NAND2X1 U6172 ( .A(n3730), .B(n1783), .Y(n4054) );
  NAND2X1 U6173 ( .A(n3730), .B(n1738), .Y(n3966) );
  NAND2X1 U6174 ( .A(n3730), .B(n1694), .Y(n3926) );
  NAND2X1 U6175 ( .A(n3730), .B(n1650), .Y(n3887) );
  NAND2X1 U6176 ( .A(n3730), .B(n1606), .Y(n3848) );
  NAND2X1 U6177 ( .A(n3730), .B(n1562), .Y(n3809) );
  NAND2X1 U6178 ( .A(n3730), .B(n1518), .Y(n3770) );
  NAND2X1 U6179 ( .A(n3730), .B(n1062), .Y(n3727) );
  NAND2X1 U6180 ( .A(n3413), .B(n1783), .Y(n3687) );
  NAND2X1 U6181 ( .A(n3413), .B(n1738), .Y(n3648) );
  NAND2X1 U6182 ( .A(n3413), .B(n1694), .Y(n3609) );
  NAND2X1 U6183 ( .A(n3413), .B(n1650), .Y(n3570) );
  NAND2X1 U6184 ( .A(n3413), .B(n1606), .Y(n3531) );
  NAND2X1 U6185 ( .A(n3413), .B(n1562), .Y(n3492) );
  NAND2X1 U6186 ( .A(n3413), .B(n1518), .Y(n3453) );
  NAND2X1 U6187 ( .A(n3413), .B(n1062), .Y(n3410) );
  NAND2X1 U6188 ( .A(n2462), .B(n1783), .Y(n2736) );
  NAND2X1 U6189 ( .A(n2462), .B(n1738), .Y(n2697) );
  NAND2X1 U6190 ( .A(n2462), .B(n1694), .Y(n2658) );
  NAND2X1 U6191 ( .A(n2462), .B(n1650), .Y(n2619) );
  NAND2X1 U6192 ( .A(n2145), .B(n1783), .Y(n2419) );
  NAND2X1 U6193 ( .A(n2145), .B(n1738), .Y(n2380) );
  NAND2X1 U6194 ( .A(n2145), .B(n1694), .Y(n2341) );
  NAND2X1 U6195 ( .A(n2145), .B(n1650), .Y(n2302) );
  NAND2X1 U6196 ( .A(n1827), .B(n1783), .Y(n2102) );
  NAND2X1 U6197 ( .A(n1827), .B(n1738), .Y(n2063) );
  NAND2X1 U6198 ( .A(n2462), .B(n1606), .Y(n2580) );
  NAND2X1 U6199 ( .A(n2462), .B(n1562), .Y(n2541) );
  NAND2X1 U6200 ( .A(n2462), .B(n1518), .Y(n2502) );
  NAND2X1 U6201 ( .A(n2462), .B(n1062), .Y(n2459) );
  NAND2X1 U6202 ( .A(n2145), .B(n1606), .Y(n2263) );
  NAND2X1 U6203 ( .A(n2145), .B(n1562), .Y(n2224) );
  NAND2X1 U6204 ( .A(n2145), .B(n1518), .Y(n2185) );
  NAND2X1 U6205 ( .A(n2145), .B(n1062), .Y(n2142) );
  NOR3X1 U6206 ( .A(n6512), .B(n6577), .C(n3364), .Y(n3359) );
  NOR3X1 U6207 ( .A(n6520), .B(n6585), .C(n3325), .Y(n3320) );
  NOR3X1 U6208 ( .A(n6528), .B(n6593), .C(n3286), .Y(n3281) );
  NOR3X1 U6209 ( .A(n6536), .B(n6601), .C(n3247), .Y(n3242) );
  NOR3X1 U6210 ( .A(n6544), .B(n6609), .C(n3208), .Y(n3203) );
  NOR3X1 U6211 ( .A(n6552), .B(n6617), .C(n3169), .Y(n3164) );
  NOR3X1 U6212 ( .A(n6560), .B(n6625), .C(n3130), .Y(n3125) );
  NOR3X1 U6213 ( .A(n6568), .B(n6633), .C(n3086), .Y(n3081) );
  NOR3X1 U6214 ( .A(n6510), .B(n6575), .C(n4047), .Y(n4042) );
  NOR3X1 U6215 ( .A(n6518), .B(n6583), .C(n3959), .Y(n3954) );
  NOR3X1 U6216 ( .A(n6526), .B(n6591), .C(n3920), .Y(n3915) );
  NOR3X1 U6217 ( .A(n6534), .B(n6599), .C(n3881), .Y(n3876) );
  NOR3X1 U6218 ( .A(n6542), .B(n6607), .C(n3842), .Y(n3837) );
  NOR3X1 U6219 ( .A(n6550), .B(n6615), .C(n3803), .Y(n3798) );
  NOR3X1 U6220 ( .A(n6558), .B(n6623), .C(n3764), .Y(n3759) );
  NOR3X1 U6221 ( .A(n6566), .B(n6631), .C(n3720), .Y(n3715) );
  NOR3X1 U6222 ( .A(n6511), .B(n6576), .C(n3681), .Y(n3676) );
  NOR3X1 U6223 ( .A(n6519), .B(n6584), .C(n3642), .Y(n3637) );
  NOR3X1 U6224 ( .A(n6527), .B(n6592), .C(n3603), .Y(n3598) );
  NOR3X1 U6225 ( .A(n6535), .B(n6600), .C(n3564), .Y(n3559) );
  NOR3X1 U6226 ( .A(n6543), .B(n6608), .C(n3525), .Y(n3520) );
  NOR3X1 U6227 ( .A(n6551), .B(n6616), .C(n3486), .Y(n3481) );
  NOR3X1 U6228 ( .A(n6559), .B(n6624), .C(n3447), .Y(n3442) );
  NOR3X1 U6229 ( .A(n6567), .B(n6632), .C(n3403), .Y(n3398) );
  NOR3X1 U6230 ( .A(n6514), .B(n6579), .C(n2730), .Y(n2725) );
  NOR3X1 U6231 ( .A(n6522), .B(n6587), .C(n2691), .Y(n2686) );
  NOR3X1 U6232 ( .A(n6530), .B(n6595), .C(n2652), .Y(n2647) );
  NOR3X1 U6233 ( .A(n6538), .B(n6603), .C(n2613), .Y(n2608) );
  NOR3X1 U6234 ( .A(n6515), .B(n6580), .C(n2413), .Y(n2408) );
  NOR3X1 U6235 ( .A(n6523), .B(n6588), .C(n2374), .Y(n2369) );
  NOR3X1 U6236 ( .A(n6531), .B(n6596), .C(n2335), .Y(n2330) );
  NOR3X1 U6237 ( .A(n6539), .B(n6604), .C(n2296), .Y(n2291) );
  NOR3X1 U6238 ( .A(n6546), .B(n6611), .C(n2574), .Y(n2569) );
  NOR3X1 U6239 ( .A(n6554), .B(n6619), .C(n2535), .Y(n2530) );
  NOR3X1 U6240 ( .A(n6562), .B(n6627), .C(n2496), .Y(n2491) );
  NOR3X1 U6241 ( .A(n6570), .B(n6635), .C(n2452), .Y(n2447) );
  NOR3X1 U6242 ( .A(n6547), .B(n6612), .C(n2257), .Y(n2252) );
  NOR3X1 U6243 ( .A(n6555), .B(n6620), .C(n2218), .Y(n2213) );
  NOR3X1 U6244 ( .A(n6563), .B(n6628), .C(n2179), .Y(n2174) );
  NOR3X1 U6245 ( .A(n6571), .B(n6636), .C(n2135), .Y(n2130) );
  AOI222X4 U6246 ( .A0(n5831), .A1(n3837), .B0(n3835), .B1(n3838), .C0(n5848), 
        .C1(n6542), .Y(n3817) );
  AO21X1 U6247 ( .A0(n5803), .A1(n6542), .B0(n3839), .Y(n3838) );
  AOI222X4 U6248 ( .A0(n5831), .A1(n3798), .B0(n3796), .B1(n3799), .C0(n5848), 
        .C1(n6550), .Y(n3778) );
  AO21X1 U6249 ( .A0(n5802), .A1(n6550), .B0(n3800), .Y(n3799) );
  AOI222X4 U6250 ( .A0(n5831), .A1(n3759), .B0(n3757), .B1(n3760), .C0(n5848), 
        .C1(n6558), .Y(n3739) );
  AO21X1 U6251 ( .A0(n5802), .A1(n6558), .B0(n3761), .Y(n3760) );
  AOI222X4 U6252 ( .A0(n5831), .A1(n3715), .B0(n3713), .B1(n3716), .C0(n5848), 
        .C1(n6566), .Y(n3695) );
  AO21X1 U6253 ( .A0(n5801), .A1(n6566), .B0(n3717), .Y(n3716) );
  AOI222X4 U6254 ( .A0(n5832), .A1(n3520), .B0(n3518), .B1(n3521), .C0(n5848), 
        .C1(n6543), .Y(n3500) );
  AO21X1 U6255 ( .A0(n5806), .A1(n6543), .B0(n3522), .Y(n3521) );
  AOI222X4 U6256 ( .A0(n5831), .A1(n3481), .B0(n3479), .B1(n3482), .C0(n5848), 
        .C1(n6551), .Y(n3461) );
  AO21X1 U6257 ( .A0(n5806), .A1(n6551), .B0(n3483), .Y(n3482) );
  AOI222X4 U6258 ( .A0(n5832), .A1(n3442), .B0(n3440), .B1(n3443), .C0(n5848), 
        .C1(n6559), .Y(n3422) );
  AO21X1 U6259 ( .A0(n5806), .A1(n6559), .B0(n3444), .Y(n3443) );
  AOI222X4 U6260 ( .A0(n5832), .A1(n3398), .B0(n3396), .B1(n3399), .C0(n5847), 
        .C1(n6567), .Y(n3378) );
  AO21X1 U6261 ( .A0(n5806), .A1(n6567), .B0(n3400), .Y(n3399) );
  AOI222X4 U6262 ( .A0(n5832), .A1(n3359), .B0(n3357), .B1(n3360), .C0(n5847), 
        .C1(n6512), .Y(n3339) );
  AO21X1 U6263 ( .A0(n5806), .A1(n6512), .B0(n3361), .Y(n3360) );
  AOI222X4 U6264 ( .A0(n5832), .A1(n3320), .B0(n3318), .B1(n3321), .C0(n5847), 
        .C1(n6520), .Y(n3300) );
  AO21X1 U6265 ( .A0(n5806), .A1(n6520), .B0(n3322), .Y(n3321) );
  AOI222X4 U6266 ( .A0(n5832), .A1(n3281), .B0(n3279), .B1(n3282), .C0(n5847), 
        .C1(n6528), .Y(n3261) );
  AO21X1 U6267 ( .A0(n5806), .A1(n6528), .B0(n3283), .Y(n3282) );
  AOI222X4 U6268 ( .A0(n5832), .A1(n3242), .B0(n3240), .B1(n3243), .C0(n5847), 
        .C1(n6536), .Y(n3222) );
  AO21X1 U6269 ( .A0(n5806), .A1(n6536), .B0(n3244), .Y(n3243) );
  AOI222X4 U6270 ( .A0(n5832), .A1(n3203), .B0(n3201), .B1(n3204), .C0(n5847), 
        .C1(n6544), .Y(n3183) );
  AO21X1 U6271 ( .A0(n5806), .A1(n6544), .B0(n3205), .Y(n3204) );
  AOI222X4 U6272 ( .A0(n5832), .A1(n3164), .B0(n3162), .B1(n3165), .C0(n5847), 
        .C1(n6552), .Y(n3144) );
  AO21X1 U6273 ( .A0(n5806), .A1(n6552), .B0(n3166), .Y(n3165) );
  AOI222X4 U6274 ( .A0(n5833), .A1(n3125), .B0(n3123), .B1(n3126), .C0(n5847), 
        .C1(n6560), .Y(n3105) );
  AO21X1 U6275 ( .A0(n5806), .A1(n6560), .B0(n3127), .Y(n3126) );
  AOI222X4 U6276 ( .A0(n5833), .A1(n3081), .B0(n3079), .B1(n3082), .C0(n5847), 
        .C1(n6568), .Y(n3061) );
  AO21X1 U6277 ( .A0(n5806), .A1(n6568), .B0(n3083), .Y(n3082) );
  AOI222X4 U6278 ( .A0(n5833), .A1(n3042), .B0(n3040), .B1(n3043), .C0(n5847), 
        .C1(n6513), .Y(n3022) );
  AO21X1 U6279 ( .A0(n5806), .A1(n6513), .B0(n3044), .Y(n3043) );
  AOI222X4 U6280 ( .A0(n5832), .A1(n3003), .B0(n3001), .B1(n3004), .C0(n5847), 
        .C1(n6521), .Y(n2983) );
  AO21X1 U6281 ( .A0(n5806), .A1(n6521), .B0(n3005), .Y(n3004) );
  AOI222X4 U6282 ( .A0(n5832), .A1(n2964), .B0(n2962), .B1(n2965), .C0(n5847), 
        .C1(n6529), .Y(n2944) );
  AO21X1 U6283 ( .A0(n5806), .A1(n6529), .B0(n2966), .Y(n2965) );
  AOI222X4 U6284 ( .A0(n5833), .A1(n2925), .B0(n2923), .B1(n2926), .C0(n5847), 
        .C1(n6537), .Y(n2905) );
  AO21X1 U6285 ( .A0(n5806), .A1(n6537), .B0(n2927), .Y(n2926) );
  AOI222X4 U6286 ( .A0(n5833), .A1(n2886), .B0(n2884), .B1(n2887), .C0(n5847), 
        .C1(n6545), .Y(n2866) );
  AO21X1 U6287 ( .A0(n5806), .A1(n6545), .B0(n2888), .Y(n2887) );
  AOI222X4 U6288 ( .A0(n5833), .A1(n2847), .B0(n2845), .B1(n2848), .C0(n5847), 
        .C1(n6553), .Y(n2827) );
  AO21X1 U6289 ( .A0(n5805), .A1(n6553), .B0(n2849), .Y(n2848) );
  AOI222X4 U6290 ( .A0(n5833), .A1(n2808), .B0(n2806), .B1(n2809), .C0(n5847), 
        .C1(n6561), .Y(n2788) );
  AO21X1 U6291 ( .A0(n5805), .A1(n6561), .B0(n2810), .Y(n2809) );
  AOI222X4 U6292 ( .A0(n5833), .A1(n2764), .B0(n2762), .B1(n2765), .C0(n5847), 
        .C1(n6569), .Y(n2744) );
  AO21X1 U6293 ( .A0(n5805), .A1(n6569), .B0(n2766), .Y(n2765) );
  AOI222X4 U6294 ( .A0(n5831), .A1(n2091), .B0(n2089), .B1(n2092), .C0(n5846), 
        .C1(n6516), .Y(n2071) );
  AO21X1 U6295 ( .A0(n5806), .A1(n6516), .B0(n2093), .Y(n2092) );
  AOI222X4 U6296 ( .A0(n5831), .A1(n2052), .B0(n2050), .B1(n2053), .C0(n5846), 
        .C1(n6524), .Y(n2032) );
  AO21X1 U6297 ( .A0(n5806), .A1(n6524), .B0(n2054), .Y(n2053) );
  AOI222X4 U6298 ( .A0(n5832), .A1(n2569), .B0(n2567), .B1(n2570), .C0(n5846), 
        .C1(n6546), .Y(n2549) );
  AO21X1 U6299 ( .A0(n5805), .A1(n6546), .B0(n2571), .Y(n2570) );
  AOI222X4 U6300 ( .A0(n5832), .A1(n2530), .B0(n2528), .B1(n2531), .C0(n5846), 
        .C1(n6554), .Y(n2510) );
  AO21X1 U6301 ( .A0(n5805), .A1(n6554), .B0(n2532), .Y(n2531) );
  AOI222X4 U6302 ( .A0(n5832), .A1(n2491), .B0(n2489), .B1(n2492), .C0(n5846), 
        .C1(n6562), .Y(n2471) );
  AO21X1 U6303 ( .A0(n5805), .A1(n6562), .B0(n2493), .Y(n2492) );
  AOI222X4 U6304 ( .A0(n5832), .A1(n2447), .B0(n2445), .B1(n2448), .C0(n5846), 
        .C1(n6570), .Y(n2427) );
  AO21X1 U6305 ( .A0(n5805), .A1(n6570), .B0(n2449), .Y(n2448) );
  AOI222X4 U6306 ( .A0(n5831), .A1(n2252), .B0(n2250), .B1(n2253), .C0(n5846), 
        .C1(n6547), .Y(n2232) );
  AO21X1 U6307 ( .A0(n5805), .A1(n6547), .B0(n2254), .Y(n2253) );
  AOI222X4 U6308 ( .A0(n5831), .A1(n2213), .B0(n2211), .B1(n2214), .C0(n5846), 
        .C1(n6555), .Y(n2193) );
  AO21X1 U6309 ( .A0(n5805), .A1(n6555), .B0(n2215), .Y(n2214) );
  AOI222X4 U6310 ( .A0(n5831), .A1(n2174), .B0(n2172), .B1(n2175), .C0(n5846), 
        .C1(n6563), .Y(n2154) );
  AO21X1 U6311 ( .A0(n5805), .A1(n6563), .B0(n2176), .Y(n2175) );
  AOI222X4 U6312 ( .A0(n5831), .A1(n2130), .B0(n2128), .B1(n2131), .C0(n5846), 
        .C1(n6571), .Y(n2110) );
  AO21X1 U6313 ( .A0(n5805), .A1(n6571), .B0(n2132), .Y(n2131) );
  OAI22X2 U6314 ( .A0(n1027), .A1(n5843), .B0(n6638), .B1(n1029), .Y(n985) );
  AOI211X1 U6315 ( .A0(n5804), .A1(n6573), .B0(n1026), .C0(n1030), .Y(n1029)
         );
  NOR3X1 U6316 ( .A(n5836), .B(n6573), .C(n1032), .Y(n1030) );
  OAI22X2 U6317 ( .A0(n5852), .A1(n1023), .B0(n1024), .B1(n1025), .Y(n986) );
  NOR2X1 U6318 ( .A(n1026), .B(n5800), .Y(n1024) );
  AOI2BB2X2 U6319 ( .B0(n5845), .B1(n6532), .A0N(n6597), .A1N(n2011), .Y(n1991) );
  AOI211X1 U6320 ( .A0(n6532), .A1(n5805), .B0(n2012), .C0(n2013), .Y(n2011)
         );
  NOR3X1 U6321 ( .A(n2014), .B(n6532), .C(n5830), .Y(n2013) );
  AOI2BB2X2 U6322 ( .B0(n5845), .B1(n6540), .A0N(n6605), .A1N(n1972), .Y(n1952) );
  AOI211X1 U6323 ( .A0(n6540), .A1(n5804), .B0(n1973), .C0(n1974), .Y(n1972)
         );
  NOR3X1 U6324 ( .A(n1975), .B(n6540), .C(n5837), .Y(n1974) );
  AOI2BB2X2 U6325 ( .B0(n5845), .B1(n6548), .A0N(n6613), .A1N(n1933), .Y(n1913) );
  AOI211X1 U6326 ( .A0(n6548), .A1(n5804), .B0(n1934), .C0(n1935), .Y(n1933)
         );
  NOR3X1 U6327 ( .A(n1936), .B(n6548), .C(n5840), .Y(n1935) );
  AOI2BB2X2 U6328 ( .B0(n5845), .B1(n6556), .A0N(n6621), .A1N(n1894), .Y(n1874) );
  AOI211X1 U6329 ( .A0(n6556), .A1(n5804), .B0(n1895), .C0(n1896), .Y(n1894)
         );
  NOR3X1 U6330 ( .A(n1897), .B(n6556), .C(n5828), .Y(n1896) );
  AOI2BB2X2 U6331 ( .B0(n5845), .B1(n6564), .A0N(n6629), .A1N(n1855), .Y(n1835) );
  AOI211X1 U6332 ( .A0(n6564), .A1(n5804), .B0(n1856), .C0(n1857), .Y(n1855)
         );
  NOR3X1 U6333 ( .A(n1858), .B(n6564), .C(n5841), .Y(n1857) );
  AOI2BB2X2 U6334 ( .B0(n5845), .B1(n6572), .A0N(n6637), .A1N(n1811), .Y(n1791) );
  AOI211X1 U6335 ( .A0(n6572), .A1(n5805), .B0(n1812), .C0(n1813), .Y(n1811)
         );
  NOR3X1 U6336 ( .A(n1814), .B(n6572), .C(n5836), .Y(n1813) );
  AOI2BB2X2 U6337 ( .B0(n5845), .B1(n6517), .A0N(n6582), .A1N(n1766), .Y(n1746) );
  AOI211X1 U6338 ( .A0(n6517), .A1(n5804), .B0(n1767), .C0(n1768), .Y(n1766)
         );
  NOR3X1 U6339 ( .A(n1769), .B(n6517), .C(n5837), .Y(n1768) );
  AOI2BB2X2 U6340 ( .B0(n5845), .B1(n6525), .A0N(n6590), .A1N(n1722), .Y(n1702) );
  AOI211X1 U6341 ( .A0(n6525), .A1(n5804), .B0(n1723), .C0(n1724), .Y(n1722)
         );
  NOR3X1 U6342 ( .A(n1725), .B(n6525), .C(n5837), .Y(n1724) );
  AOI2BB2X2 U6343 ( .B0(n5845), .B1(n6533), .A0N(n6598), .A1N(n1678), .Y(n1658) );
  AOI211X1 U6344 ( .A0(n6533), .A1(n5804), .B0(n1679), .C0(n1680), .Y(n1678)
         );
  NOR3X1 U6345 ( .A(n1681), .B(n6533), .C(n5837), .Y(n1680) );
  AOI2BB2X2 U6346 ( .B0(n5845), .B1(n6541), .A0N(n6606), .A1N(n1634), .Y(n1614) );
  AOI211X1 U6347 ( .A0(n6541), .A1(n5804), .B0(n1635), .C0(n1636), .Y(n1634)
         );
  NOR3X1 U6348 ( .A(n1637), .B(n6541), .C(n5837), .Y(n1636) );
  AOI2BB2X2 U6349 ( .B0(n5845), .B1(n6549), .A0N(n6614), .A1N(n1590), .Y(n1570) );
  AOI211X1 U6350 ( .A0(n6549), .A1(n5804), .B0(n1591), .C0(n1592), .Y(n1590)
         );
  NOR3X1 U6351 ( .A(n1593), .B(n6549), .C(n5837), .Y(n1592) );
  AOI2BB2X2 U6352 ( .B0(n5845), .B1(n6557), .A0N(n6622), .A1N(n1546), .Y(n1526) );
  AOI211X1 U6353 ( .A0(n6557), .A1(n5804), .B0(n1547), .C0(n1548), .Y(n1546)
         );
  NOR3X1 U6354 ( .A(n1549), .B(n6557), .C(n5837), .Y(n1548) );
  AOI2BB2X2 U6355 ( .B0(n5845), .B1(n6565), .A0N(n6630), .A1N(n1502), .Y(n1482) );
  AOI211X1 U6356 ( .A0(n6565), .A1(n5804), .B0(n1503), .C0(n1504), .Y(n1502)
         );
  NOR3X1 U6357 ( .A(n1505), .B(n6565), .C(n5836), .Y(n1504) );
  INVX3 U6358 ( .A(n1585), .Y(n6494) );
  OAI222XL U6359 ( .A0(n5814), .A1(n1586), .B0(n1587), .B1(n1588), .C0(n5815), 
        .C1(n1589), .Y(n1585) );
  OA21XL U6360 ( .A0(n6549), .A1(n5850), .B0(n5828), .Y(n1587) );
  INVX3 U6361 ( .A(n1541), .Y(n6496) );
  OAI222XL U6362 ( .A0(n5814), .A1(n1542), .B0(n1543), .B1(n1544), .C0(n5821), 
        .C1(n1545), .Y(n1541) );
  OA21XL U6363 ( .A0(n6557), .A1(n5849), .B0(n5837), .Y(n1543) );
  INVX3 U6364 ( .A(n1497), .Y(n6498) );
  OAI222XL U6365 ( .A0(n5814), .A1(n1498), .B0(n1499), .B1(n1500), .C0(n5820), 
        .C1(n1501), .Y(n1497) );
  OA21XL U6366 ( .A0(n6565), .A1(n5849), .B0(n5837), .Y(n1499) );
  OA22X2 U6367 ( .A0(n5854), .A1(n4038), .B0(n4045), .B1(n4040), .Y(n3987) );
  NOR2X1 U6368 ( .A(n4044), .B(n5799), .Y(n4045) );
  OA22X2 U6369 ( .A0(n5853), .A1(n2721), .B0(n2728), .B1(n2723), .Y(n2704) );
  NOR2X1 U6370 ( .A(n2727), .B(n5803), .Y(n2728) );
  OA22X2 U6371 ( .A0(n5853), .A1(n2682), .B0(n2689), .B1(n2684), .Y(n2665) );
  NOR2X1 U6372 ( .A(n2688), .B(n5803), .Y(n2689) );
  OA22X2 U6373 ( .A0(n5853), .A1(n2643), .B0(n2650), .B1(n2645), .Y(n2626) );
  NOR2X1 U6374 ( .A(n2649), .B(n5803), .Y(n2650) );
  OA22X2 U6375 ( .A0(n5853), .A1(n2604), .B0(n2611), .B1(n2606), .Y(n2587) );
  NOR2X1 U6376 ( .A(n2610), .B(n5803), .Y(n2611) );
  OA22X2 U6377 ( .A0(n5853), .A1(n2404), .B0(n2411), .B1(n2406), .Y(n2387) );
  NOR2X1 U6378 ( .A(n2410), .B(n5804), .Y(n2411) );
  OA22X2 U6379 ( .A0(n5853), .A1(n2365), .B0(n2372), .B1(n2367), .Y(n2348) );
  NOR2X1 U6380 ( .A(n2371), .B(n5803), .Y(n2372) );
  OA22X2 U6381 ( .A0(n5853), .A1(n2326), .B0(n2333), .B1(n2328), .Y(n2309) );
  NOR2X1 U6382 ( .A(n2332), .B(n5803), .Y(n2333) );
  OA22X2 U6383 ( .A0(n5853), .A1(n2287), .B0(n2294), .B1(n2289), .Y(n2270) );
  NOR2X1 U6384 ( .A(n2293), .B(n5803), .Y(n2294) );
  OA22X2 U6385 ( .A0(n5852), .A1(n2007), .B0(n2015), .B1(n2009), .Y(n1990) );
  NOR2X1 U6386 ( .A(n2012), .B(n5802), .Y(n2015) );
  OA22X2 U6387 ( .A0(n5852), .A1(n1968), .B0(n1976), .B1(n1970), .Y(n1951) );
  NOR2X1 U6388 ( .A(n1973), .B(n5802), .Y(n1976) );
  OA22X2 U6389 ( .A0(n5852), .A1(n1929), .B0(n1937), .B1(n1931), .Y(n1912) );
  NOR2X1 U6390 ( .A(n1934), .B(n5801), .Y(n1937) );
  OA22X2 U6391 ( .A0(n5852), .A1(n1890), .B0(n1898), .B1(n1892), .Y(n1873) );
  NOR2X1 U6392 ( .A(n1895), .B(n5801), .Y(n1898) );
  OA22X2 U6393 ( .A0(n5852), .A1(n1851), .B0(n1859), .B1(n1853), .Y(n1834) );
  NOR2X1 U6394 ( .A(n1856), .B(n5801), .Y(n1859) );
  OA22X2 U6395 ( .A0(n5852), .A1(n1807), .B0(n1815), .B1(n1809), .Y(n1790) );
  NOR2X1 U6396 ( .A(n1812), .B(n5801), .Y(n1815) );
  OA22X2 U6397 ( .A0(n5852), .A1(n1762), .B0(n1770), .B1(n1764), .Y(n1745) );
  NOR2X1 U6398 ( .A(n1767), .B(n5800), .Y(n1770) );
  OA22X2 U6399 ( .A0(n5852), .A1(n1718), .B0(n1726), .B1(n1720), .Y(n1701) );
  NOR2X1 U6400 ( .A(n1723), .B(n5800), .Y(n1726) );
  OA22X2 U6401 ( .A0(n5852), .A1(n1674), .B0(n1682), .B1(n1676), .Y(n1657) );
  NOR2X1 U6402 ( .A(n1679), .B(n5800), .Y(n1682) );
  OA22X2 U6403 ( .A0(n5852), .A1(n1630), .B0(n1638), .B1(n1632), .Y(n1613) );
  NOR2X1 U6404 ( .A(n1635), .B(n5800), .Y(n1638) );
  OA22X2 U6405 ( .A0(n5852), .A1(n1586), .B0(n1594), .B1(n1588), .Y(n1569) );
  NOR2X1 U6406 ( .A(n1591), .B(n5799), .Y(n1594) );
  OA22X2 U6407 ( .A0(n5852), .A1(n1542), .B0(n1550), .B1(n1544), .Y(n1525) );
  NOR2X1 U6408 ( .A(n1547), .B(n5799), .Y(n1550) );
  OA22X2 U6409 ( .A0(n5852), .A1(n1498), .B0(n1506), .B1(n1500), .Y(n1481) );
  NOR2X1 U6410 ( .A(n1503), .B(n5799), .Y(n1506) );
  AO22X2 U6411 ( .A0(n4042), .A1(n5764), .B0(n6510), .B1(n4046), .Y(n3971) );
  AO22X1 U6412 ( .A0(n4040), .A1(n5833), .B0(n4041), .B1(n5823), .Y(n4046) );
  AO22X2 U6413 ( .A0(n3954), .A1(n5764), .B0(n6518), .B1(n3958), .Y(n3931) );
  AO22X1 U6414 ( .A0(n3952), .A1(n5834), .B0(n3953), .B1(n5822), .Y(n3958) );
  AO22X2 U6415 ( .A0(n3915), .A1(n5764), .B0(n6526), .B1(n3919), .Y(n3892) );
  AO22X1 U6416 ( .A0(n3913), .A1(n5834), .B0(n3914), .B1(n5825), .Y(n3919) );
  AO22X2 U6417 ( .A0(n3876), .A1(n5764), .B0(n6534), .B1(n3880), .Y(n3853) );
  AO22X1 U6418 ( .A0(n3874), .A1(n5832), .B0(n3875), .B1(n5822), .Y(n3880) );
  AO22X2 U6419 ( .A0(n3837), .A1(n5764), .B0(n6542), .B1(n3841), .Y(n3814) );
  AO22X1 U6420 ( .A0(n3835), .A1(n5834), .B0(n3836), .B1(n5824), .Y(n3841) );
  AO22X2 U6421 ( .A0(n3798), .A1(n5764), .B0(n6550), .B1(n3802), .Y(n3775) );
  AO22X1 U6422 ( .A0(n3796), .A1(n5832), .B0(n3797), .B1(n5823), .Y(n3802) );
  AO22X2 U6423 ( .A0(n3759), .A1(n5764), .B0(n6558), .B1(n3763), .Y(n3736) );
  AO22X1 U6424 ( .A0(n3757), .A1(n5832), .B0(n3758), .B1(n5822), .Y(n3763) );
  AO22X2 U6425 ( .A0(n3715), .A1(n5764), .B0(n6566), .B1(n3719), .Y(n3692) );
  AO22X1 U6426 ( .A0(n3713), .A1(n5832), .B0(n3714), .B1(n5823), .Y(n3719) );
  AO22X2 U6427 ( .A0(n3676), .A1(n5764), .B0(n6511), .B1(n3680), .Y(n3653) );
  AO22X1 U6428 ( .A0(n3674), .A1(n5832), .B0(n3675), .B1(n5822), .Y(n3680) );
  AO22X2 U6429 ( .A0(n3637), .A1(n5764), .B0(n6519), .B1(n3641), .Y(n3614) );
  AO22X1 U6430 ( .A0(n3635), .A1(n5834), .B0(n3636), .B1(n5825), .Y(n3641) );
  AO22X2 U6431 ( .A0(n3598), .A1(n5764), .B0(n6527), .B1(n3602), .Y(n3575) );
  AO22X1 U6432 ( .A0(n3596), .A1(n5832), .B0(n3597), .B1(n5823), .Y(n3602) );
  AO22X2 U6433 ( .A0(n3559), .A1(n5764), .B0(n6535), .B1(n3563), .Y(n3536) );
  AO22X1 U6434 ( .A0(n3557), .A1(n5834), .B0(n3558), .B1(n5825), .Y(n3563) );
  AO22X2 U6435 ( .A0(n3520), .A1(n5764), .B0(n6543), .B1(n3524), .Y(n3497) );
  AO22X1 U6436 ( .A0(n3518), .A1(n5834), .B0(n3519), .B1(n5823), .Y(n3524) );
  AO22X2 U6437 ( .A0(n3481), .A1(n5764), .B0(n6551), .B1(n3485), .Y(n3458) );
  AO22X1 U6438 ( .A0(n3479), .A1(n5834), .B0(n3480), .B1(n5822), .Y(n3485) );
  AO22X2 U6439 ( .A0(n3442), .A1(n5764), .B0(n6559), .B1(n3446), .Y(n3419) );
  AO22X1 U6440 ( .A0(n3440), .A1(n5834), .B0(n3441), .B1(n5822), .Y(n3446) );
  AO22X2 U6441 ( .A0(n3398), .A1(n5764), .B0(n6567), .B1(n3402), .Y(n3375) );
  AO22X1 U6442 ( .A0(n3396), .A1(n5834), .B0(n3397), .B1(n5827), .Y(n3402) );
  AO22X2 U6443 ( .A0(n3359), .A1(n5764), .B0(n6512), .B1(n3363), .Y(n3336) );
  AO22X1 U6444 ( .A0(n3357), .A1(n5834), .B0(n3358), .B1(n5827), .Y(n3363) );
  AO22X2 U6445 ( .A0(n3320), .A1(n5764), .B0(n6520), .B1(n3324), .Y(n3297) );
  AO22X1 U6446 ( .A0(n3318), .A1(n5834), .B0(n3319), .B1(n5827), .Y(n3324) );
  AO22X2 U6447 ( .A0(n3281), .A1(n5764), .B0(n6528), .B1(n3285), .Y(n3258) );
  AO22X1 U6448 ( .A0(n3279), .A1(n5834), .B0(n3280), .B1(n5823), .Y(n3285) );
  AO22X2 U6449 ( .A0(n3242), .A1(n5764), .B0(n6536), .B1(n3246), .Y(n3219) );
  AO22X1 U6450 ( .A0(n3240), .A1(n5834), .B0(n3241), .B1(n5823), .Y(n3246) );
  AO22X2 U6451 ( .A0(n3203), .A1(n5764), .B0(n6544), .B1(n3207), .Y(n3180) );
  AO22X1 U6452 ( .A0(n3201), .A1(n5834), .B0(n3202), .B1(n5824), .Y(n3207) );
  AO22X2 U6453 ( .A0(n3164), .A1(n5764), .B0(n6552), .B1(n3168), .Y(n3141) );
  AO22X1 U6454 ( .A0(n3162), .A1(n5834), .B0(n3163), .B1(n5822), .Y(n3168) );
  AO22X2 U6455 ( .A0(n3125), .A1(n5764), .B0(n6560), .B1(n3129), .Y(n3102) );
  AO22X1 U6456 ( .A0(n3123), .A1(n5834), .B0(n3124), .B1(n5822), .Y(n3129) );
  AO22X2 U6457 ( .A0(n3081), .A1(n5765), .B0(n6568), .B1(n3085), .Y(n3058) );
  AO22X1 U6458 ( .A0(n3079), .A1(n5834), .B0(n3080), .B1(n5824), .Y(n3085) );
  AO22X2 U6459 ( .A0(n3042), .A1(n5765), .B0(n6513), .B1(n3046), .Y(n3019) );
  AO22X1 U6460 ( .A0(n3040), .A1(n5834), .B0(n3041), .B1(n5824), .Y(n3046) );
  AO22X2 U6461 ( .A0(n3003), .A1(n5765), .B0(n6521), .B1(n3007), .Y(n2980) );
  AO22X1 U6462 ( .A0(n3001), .A1(n5834), .B0(n3002), .B1(n5822), .Y(n3007) );
  AO22X2 U6463 ( .A0(n2964), .A1(n5765), .B0(n6529), .B1(n2968), .Y(n2941) );
  AO22X1 U6464 ( .A0(n2962), .A1(n5834), .B0(n2963), .B1(n5822), .Y(n2968) );
  AO22X2 U6465 ( .A0(n2925), .A1(n5765), .B0(n6537), .B1(n2929), .Y(n2902) );
  AO22X1 U6466 ( .A0(n2923), .A1(n5834), .B0(n2924), .B1(n5825), .Y(n2929) );
  AO22X2 U6467 ( .A0(n2886), .A1(n5765), .B0(n6545), .B1(n2890), .Y(n2863) );
  AO22X1 U6468 ( .A0(n2884), .A1(n5834), .B0(n2885), .B1(n5824), .Y(n2890) );
  AO22X2 U6469 ( .A0(n2847), .A1(n5765), .B0(n6553), .B1(n2851), .Y(n2824) );
  AO22X1 U6470 ( .A0(n2845), .A1(n5834), .B0(n2846), .B1(n5822), .Y(n2851) );
  AO22X2 U6471 ( .A0(n2808), .A1(n5765), .B0(n6561), .B1(n2812), .Y(n2785) );
  AO22X1 U6472 ( .A0(n2806), .A1(n5834), .B0(n2807), .B1(n5824), .Y(n2812) );
  AO22X2 U6473 ( .A0(n2764), .A1(n5765), .B0(n6569), .B1(n2768), .Y(n2741) );
  AO22X1 U6474 ( .A0(n2762), .A1(n5834), .B0(n2763), .B1(n5823), .Y(n2768) );
  AO22X2 U6475 ( .A0(n2725), .A1(n5765), .B0(n6514), .B1(n2729), .Y(n2702) );
  AO22X1 U6476 ( .A0(n2723), .A1(n5834), .B0(n2724), .B1(n5822), .Y(n2729) );
  AO22X2 U6477 ( .A0(n2686), .A1(n5765), .B0(n6522), .B1(n2690), .Y(n2663) );
  AO22X1 U6478 ( .A0(n2684), .A1(n5834), .B0(n2685), .B1(n5822), .Y(n2690) );
  AO22X2 U6479 ( .A0(n2647), .A1(n5765), .B0(n6530), .B1(n2651), .Y(n2624) );
  AO22X1 U6480 ( .A0(n2645), .A1(n5834), .B0(n2646), .B1(n5825), .Y(n2651) );
  AO22X2 U6481 ( .A0(n2608), .A1(n5765), .B0(n6538), .B1(n2612), .Y(n2585) );
  AO22X1 U6482 ( .A0(n2606), .A1(n5833), .B0(n2607), .B1(n5824), .Y(n2612) );
  AO22X2 U6483 ( .A0(n2569), .A1(n5765), .B0(n6546), .B1(n2573), .Y(n2546) );
  AO22X1 U6484 ( .A0(n2567), .A1(n5833), .B0(n2568), .B1(n5823), .Y(n2573) );
  AO22X2 U6485 ( .A0(n2530), .A1(n5765), .B0(n6554), .B1(n2534), .Y(n2507) );
  AO22X1 U6486 ( .A0(n2528), .A1(n5833), .B0(n2529), .B1(n5823), .Y(n2534) );
  AO22X2 U6487 ( .A0(n2491), .A1(n5765), .B0(n6562), .B1(n2495), .Y(n2468) );
  AO22X1 U6488 ( .A0(n2489), .A1(n5833), .B0(n2490), .B1(n5823), .Y(n2495) );
  AO22X2 U6489 ( .A0(n2447), .A1(n5765), .B0(n6570), .B1(n2451), .Y(n2424) );
  AO22X1 U6490 ( .A0(n2445), .A1(n5833), .B0(n2446), .B1(n5822), .Y(n2451) );
  AO22X2 U6491 ( .A0(n2408), .A1(n5765), .B0(n6515), .B1(n2412), .Y(n2385) );
  AO22X1 U6492 ( .A0(n2406), .A1(n5833), .B0(n2407), .B1(n5827), .Y(n2412) );
  AO22X2 U6493 ( .A0(n2369), .A1(n5765), .B0(n6523), .B1(n2373), .Y(n2346) );
  AO22X1 U6494 ( .A0(n2367), .A1(n5834), .B0(n2368), .B1(n5823), .Y(n2373) );
  AO22X2 U6495 ( .A0(n2330), .A1(n5765), .B0(n6531), .B1(n2334), .Y(n2307) );
  AO22X1 U6496 ( .A0(n2328), .A1(n5833), .B0(n2329), .B1(n5823), .Y(n2334) );
  AO22X2 U6497 ( .A0(n2291), .A1(n5765), .B0(n6539), .B1(n2295), .Y(n2268) );
  AO22X1 U6498 ( .A0(n2289), .A1(n5833), .B0(n2290), .B1(n5822), .Y(n2295) );
  AO22X2 U6499 ( .A0(n2252), .A1(n5765), .B0(n6547), .B1(n2256), .Y(n2229) );
  AO22X1 U6500 ( .A0(n2250), .A1(n5833), .B0(n2251), .B1(n5824), .Y(n2256) );
  AO22X2 U6501 ( .A0(n2213), .A1(n5765), .B0(n6555), .B1(n2217), .Y(n2190) );
  AO22X1 U6502 ( .A0(n2211), .A1(n5833), .B0(n2212), .B1(n5824), .Y(n2217) );
  AO22X2 U6503 ( .A0(n2174), .A1(n5765), .B0(n6563), .B1(n2178), .Y(n2151) );
  AO22X1 U6504 ( .A0(n2172), .A1(n5833), .B0(n2173), .B1(n5824), .Y(n2178) );
  AO22X2 U6505 ( .A0(n2130), .A1(n5765), .B0(n6571), .B1(n2134), .Y(n2107) );
  AO22X1 U6506 ( .A0(n2128), .A1(n5833), .B0(n2129), .B1(n5823), .Y(n2134) );
  INVX3 U6507 ( .A(n1640), .Y(n6491) );
  AOI32X1 U6508 ( .A0(n6541), .A1(n1633), .A2(n5825), .B0(n1632), .B1(n1641), 
        .Y(n1640) );
  OAI32X1 U6509 ( .A0(n4827), .A1(n6541), .A2(n1637), .B0(n1639), .B1(n5835), 
        .Y(n1641) );
  AOI32X4 U6510 ( .A0(n5824), .A1(n1033), .A2(n6573), .B0(n1025), .B1(n1038), 
        .Y(n982) );
  OAI32X1 U6511 ( .A0(n4827), .A1(n6573), .A2(n1032), .B0(n5838), .B1(n1027), 
        .Y(n1038) );
  INVX3 U6512 ( .A(n1552), .Y(n6495) );
  AOI32X1 U6513 ( .A0(n6557), .A1(n1545), .A2(n5825), .B0(n1544), .B1(n1553), 
        .Y(n1552) );
  OAI32X1 U6514 ( .A0(n4827), .A1(n6557), .A2(n1549), .B0(n1551), .B1(n5838), 
        .Y(n1553) );
  INVX3 U6515 ( .A(n1508), .Y(n6497) );
  AOI32X1 U6516 ( .A0(n6565), .A1(n1501), .A2(n5825), .B0(n1500), .B1(n1509), 
        .Y(n1508) );
  OAI32X1 U6517 ( .A0(n4827), .A1(n6565), .A2(n1505), .B0(n1507), .B1(n5838), 
        .Y(n1509) );
  NAND2X1 U6518 ( .A(n1783), .B(n1061), .Y(n1771) );
  NAND2X1 U6519 ( .A(n1738), .B(n1061), .Y(n1727) );
  NAND2X1 U6520 ( .A(n1694), .B(n1061), .Y(n1683) );
  NAND2X1 U6521 ( .A(n1650), .B(n1061), .Y(n1639) );
  NAND2X1 U6522 ( .A(n1606), .B(n1061), .Y(n1595) );
  NAND2X1 U6523 ( .A(n1562), .B(n1061), .Y(n1551) );
  NAND2X1 U6524 ( .A(n1518), .B(n1061), .Y(n1507) );
  NAND2X1 U6525 ( .A(n1827), .B(n1694), .Y(n2016) );
  NAND2X1 U6526 ( .A(n1827), .B(n1650), .Y(n1977) );
  NAND2X1 U6527 ( .A(n1827), .B(n1606), .Y(n1938) );
  NAND2X1 U6528 ( .A(n1827), .B(n1562), .Y(n1899) );
  NAND2X1 U6529 ( .A(n1827), .B(n1518), .Y(n1860) );
  NAND2X1 U6530 ( .A(n1827), .B(n1062), .Y(n1816) );
  INVX3 U6531 ( .A(n4037), .Y(n6423) );
  OAI222XL U6532 ( .A0(n5813), .A1(n4038), .B0(n4039), .B1(n4040), .C0(n5821), 
        .C1(n4041), .Y(n4037) );
  OA21XL U6533 ( .A0(n6510), .A1(n5849), .B0(n5836), .Y(n4039) );
  INVX3 U6534 ( .A(n2720), .Y(n6455) );
  OAI222XL U6535 ( .A0(n5812), .A1(n2721), .B0(n2722), .B1(n2723), .C0(n5821), 
        .C1(n2724), .Y(n2720) );
  OA21XL U6536 ( .A0(n6514), .A1(n5849), .B0(n5837), .Y(n2722) );
  INVX3 U6537 ( .A(n2681), .Y(n6456) );
  OAI222XL U6538 ( .A0(n5811), .A1(n2682), .B0(n2683), .B1(n2684), .C0(n5820), 
        .C1(n2685), .Y(n2681) );
  OA21XL U6539 ( .A0(n6522), .A1(n5843), .B0(n5830), .Y(n2683) );
  INVX3 U6540 ( .A(n2642), .Y(n6457) );
  OAI222XL U6541 ( .A0(n5811), .A1(n2643), .B0(n2644), .B1(n2645), .C0(n5820), 
        .C1(n2646), .Y(n2642) );
  OA21XL U6542 ( .A0(n6530), .A1(n5849), .B0(n5839), .Y(n2644) );
  INVX3 U6543 ( .A(n2603), .Y(n6458) );
  OAI222XL U6544 ( .A0(n5814), .A1(n2604), .B0(n2605), .B1(n2606), .C0(n5820), 
        .C1(n2607), .Y(n2603) );
  OA21XL U6545 ( .A0(n6538), .A1(n5849), .B0(n5840), .Y(n2605) );
  INVX3 U6546 ( .A(n2403), .Y(n6463) );
  OAI222XL U6547 ( .A0(n5814), .A1(n2404), .B0(n2405), .B1(n2406), .C0(n5821), 
        .C1(n2407), .Y(n2403) );
  OA21XL U6548 ( .A0(n6515), .A1(n5850), .B0(n5840), .Y(n2405) );
  INVX3 U6549 ( .A(n2364), .Y(n6464) );
  OAI222XL U6550 ( .A0(n5813), .A1(n2365), .B0(n2366), .B1(n2367), .C0(n5821), 
        .C1(n2368), .Y(n2364) );
  OA21XL U6551 ( .A0(n6523), .A1(n5850), .B0(n5840), .Y(n2366) );
  INVX3 U6552 ( .A(n2325), .Y(n6465) );
  OAI222XL U6553 ( .A0(n5811), .A1(n2326), .B0(n2327), .B1(n2328), .C0(n5821), 
        .C1(n2329), .Y(n2325) );
  OA21XL U6554 ( .A0(n6531), .A1(n5850), .B0(n5828), .Y(n2327) );
  INVX3 U6555 ( .A(n2286), .Y(n6466) );
  OAI222XL U6556 ( .A0(n5813), .A1(n2287), .B0(n2288), .B1(n2289), .C0(n5821), 
        .C1(n2290), .Y(n2286) );
  OA21XL U6557 ( .A0(n6539), .A1(n5850), .B0(n5828), .Y(n2288) );
  INVX3 U6558 ( .A(n1761), .Y(n6486) );
  OAI222XL U6559 ( .A0(n5814), .A1(n1762), .B0(n1763), .B1(n1764), .C0(n5819), 
        .C1(n1765), .Y(n1761) );
  OA21XL U6560 ( .A0(n6517), .A1(n5850), .B0(n5839), .Y(n1763) );
  INVX3 U6561 ( .A(n1717), .Y(n6488) );
  OAI222XL U6562 ( .A0(n5814), .A1(n1718), .B0(n1719), .B1(n1720), .C0(n5816), 
        .C1(n1721), .Y(n1717) );
  OA21XL U6563 ( .A0(n6525), .A1(n5844), .B0(n5839), .Y(n1719) );
  INVX3 U6564 ( .A(n1673), .Y(n6490) );
  OAI222XL U6565 ( .A0(n5814), .A1(n1674), .B0(n1675), .B1(n1676), .C0(n5820), 
        .C1(n1677), .Y(n1673) );
  OA21XL U6566 ( .A0(n6533), .A1(n5849), .B0(n5839), .Y(n1675) );
  INVX3 U6567 ( .A(n1629), .Y(n6492) );
  OAI222XL U6568 ( .A0(n5814), .A1(n1630), .B0(n1631), .B1(n1632), .C0(n5820), 
        .C1(n1633), .Y(n1629) );
  OA21XL U6569 ( .A0(n6541), .A1(n5849), .B0(n5837), .Y(n1631) );
  INVX3 U6570 ( .A(n2017), .Y(n6473) );
  AOI32X1 U6571 ( .A0(n6532), .A1(n2010), .A2(n5825), .B0(n2009), .B1(n2018), 
        .Y(n2017) );
  OAI32X1 U6572 ( .A0(n4827), .A1(n6532), .A2(n2014), .B0(n2016), .B1(n5838), 
        .Y(n2018) );
  INVX3 U6573 ( .A(n1978), .Y(n6475) );
  AOI32X1 U6574 ( .A0(n6540), .A1(n1971), .A2(n5823), .B0(n1970), .B1(n1979), 
        .Y(n1978) );
  OAI32X1 U6575 ( .A0(n4827), .A1(n6540), .A2(n1975), .B0(n1977), .B1(n5842), 
        .Y(n1979) );
  INVX3 U6576 ( .A(n1939), .Y(n6477) );
  AOI32X1 U6577 ( .A0(n6548), .A1(n1932), .A2(n5824), .B0(n1931), .B1(n1940), 
        .Y(n1939) );
  OAI32X1 U6578 ( .A0(n5766), .A1(n6548), .A2(n1936), .B0(n1938), .B1(n5838), 
        .Y(n1940) );
  INVX3 U6579 ( .A(n1900), .Y(n6479) );
  AOI32X1 U6580 ( .A0(n6556), .A1(n1893), .A2(n5825), .B0(n1892), .B1(n1901), 
        .Y(n1900) );
  OAI32X1 U6581 ( .A0(n4827), .A1(n6556), .A2(n1897), .B0(n1899), .B1(n5838), 
        .Y(n1901) );
  INVX3 U6582 ( .A(n1861), .Y(n6481) );
  AOI32X1 U6583 ( .A0(n6564), .A1(n1854), .A2(n5826), .B0(n1853), .B1(n1862), 
        .Y(n1861) );
  OAI32X1 U6584 ( .A0(n4827), .A1(n6564), .A2(n1858), .B0(n1860), .B1(n5838), 
        .Y(n1862) );
  INVX3 U6585 ( .A(n1817), .Y(n6483) );
  AOI32X1 U6586 ( .A0(n6572), .A1(n1810), .A2(n5824), .B0(n1809), .B1(n1818), 
        .Y(n1817) );
  OAI32X1 U6587 ( .A0(n4827), .A1(n6572), .A2(n1814), .B0(n1816), .B1(n5838), 
        .Y(n1818) );
  INVX3 U6588 ( .A(n1772), .Y(n6485) );
  AOI32X1 U6589 ( .A0(n6517), .A1(n1765), .A2(n5825), .B0(n1764), .B1(n1773), 
        .Y(n1772) );
  OAI32X1 U6590 ( .A0(n4827), .A1(n6517), .A2(n1769), .B0(n1771), .B1(n5838), 
        .Y(n1773) );
  INVX3 U6591 ( .A(n1728), .Y(n6487) );
  AOI32X1 U6592 ( .A0(n6525), .A1(n1721), .A2(n5824), .B0(n1720), .B1(n1729), 
        .Y(n1728) );
  OAI32X1 U6593 ( .A0(n5766), .A1(n6525), .A2(n1725), .B0(n1727), .B1(n5838), 
        .Y(n1729) );
  INVX3 U6594 ( .A(n1684), .Y(n6489) );
  AOI32X1 U6595 ( .A0(n6533), .A1(n1677), .A2(n5825), .B0(n1676), .B1(n1685), 
        .Y(n1684) );
  OAI32X1 U6596 ( .A0(n5766), .A1(n6533), .A2(n1681), .B0(n1683), .B1(n5839), 
        .Y(n1685) );
  INVX3 U6597 ( .A(n1596), .Y(n6493) );
  AOI32X1 U6598 ( .A0(n6549), .A1(n1589), .A2(n5826), .B0(n1588), .B1(n1597), 
        .Y(n1596) );
  OAI32X1 U6599 ( .A0(n4827), .A1(n6549), .A2(n1593), .B0(n1595), .B1(n5838), 
        .Y(n1597) );
  NAND3X1 U6600 ( .A(n1025), .B(n1032), .C(n1027), .Y(n1023) );
  NOR3X1 U6601 ( .A(n6513), .B(n6578), .C(n3047), .Y(n3042) );
  NOR3X1 U6602 ( .A(n6521), .B(n6586), .C(n3008), .Y(n3003) );
  NOR3X1 U6603 ( .A(n6529), .B(n6594), .C(n2969), .Y(n2964) );
  NOR3X1 U6604 ( .A(n6537), .B(n6602), .C(n2930), .Y(n2925) );
  NOR3X1 U6605 ( .A(n6545), .B(n6610), .C(n2891), .Y(n2886) );
  NOR3X1 U6606 ( .A(n6553), .B(n6618), .C(n2852), .Y(n2847) );
  NOR3X1 U6607 ( .A(n6561), .B(n6626), .C(n2813), .Y(n2808) );
  NOR3X1 U6608 ( .A(n6569), .B(n6634), .C(n2769), .Y(n2764) );
  NOR3X1 U6609 ( .A(n6516), .B(n6581), .C(n2096), .Y(n2091) );
  NOR3X1 U6610 ( .A(n6524), .B(n6589), .C(n2057), .Y(n2052) );
  NAND3X1 U6611 ( .A(n4040), .B(n4047), .C(n4054), .Y(n4038) );
  NAND3X1 U6612 ( .A(n3952), .B(n3959), .C(n3966), .Y(n3950) );
  NAND3X1 U6613 ( .A(n3913), .B(n3920), .C(n3926), .Y(n3911) );
  NAND3X1 U6614 ( .A(n3874), .B(n3881), .C(n3887), .Y(n3872) );
  NAND3X1 U6615 ( .A(n3674), .B(n3681), .C(n3687), .Y(n3672) );
  NAND3X1 U6616 ( .A(n3635), .B(n3642), .C(n3648), .Y(n3633) );
  NAND3X1 U6617 ( .A(n3596), .B(n3603), .C(n3609), .Y(n3594) );
  NAND3X1 U6618 ( .A(n3557), .B(n3564), .C(n3570), .Y(n3555) );
  NAND3X1 U6619 ( .A(n3357), .B(n3364), .C(n3370), .Y(n3355) );
  NAND3X1 U6620 ( .A(n3318), .B(n3325), .C(n3331), .Y(n3316) );
  NAND3X1 U6621 ( .A(n3279), .B(n3286), .C(n3292), .Y(n3277) );
  NAND3X1 U6622 ( .A(n3240), .B(n3247), .C(n3253), .Y(n3238) );
  NAND3X1 U6623 ( .A(n3040), .B(n3047), .C(n3053), .Y(n3038) );
  NAND3X1 U6624 ( .A(n3001), .B(n3008), .C(n3014), .Y(n2999) );
  NAND3X1 U6625 ( .A(n2962), .B(n2969), .C(n2975), .Y(n2960) );
  NAND3X1 U6626 ( .A(n2923), .B(n2930), .C(n2936), .Y(n2921) );
  NAND3X1 U6627 ( .A(n2723), .B(n2730), .C(n2736), .Y(n2721) );
  NAND3X1 U6628 ( .A(n2684), .B(n2691), .C(n2697), .Y(n2682) );
  NAND3X1 U6629 ( .A(n2645), .B(n2652), .C(n2658), .Y(n2643) );
  NAND3X1 U6630 ( .A(n2606), .B(n2613), .C(n2619), .Y(n2604) );
  NAND3X1 U6631 ( .A(n2406), .B(n2413), .C(n2419), .Y(n2404) );
  NAND3X1 U6632 ( .A(n2367), .B(n2374), .C(n2380), .Y(n2365) );
  NAND3X1 U6633 ( .A(n2328), .B(n2335), .C(n2341), .Y(n2326) );
  NAND3X1 U6634 ( .A(n2289), .B(n2296), .C(n2302), .Y(n2287) );
  NAND3X1 U6635 ( .A(n2089), .B(n2096), .C(n2102), .Y(n2087) );
  NAND3X1 U6636 ( .A(n2050), .B(n2057), .C(n2063), .Y(n2048) );
  NAND3X1 U6637 ( .A(n3835), .B(n3842), .C(n3848), .Y(n3833) );
  NAND3X1 U6638 ( .A(n3796), .B(n3803), .C(n3809), .Y(n3794) );
  NAND3X1 U6639 ( .A(n3757), .B(n3764), .C(n3770), .Y(n3755) );
  NAND3X1 U6640 ( .A(n3713), .B(n3720), .C(n3727), .Y(n3711) );
  NAND3X1 U6641 ( .A(n3518), .B(n3525), .C(n3531), .Y(n3516) );
  NAND3X1 U6642 ( .A(n3479), .B(n3486), .C(n3492), .Y(n3477) );
  NAND3X1 U6643 ( .A(n3440), .B(n3447), .C(n3453), .Y(n3438) );
  NAND3X1 U6644 ( .A(n3396), .B(n3403), .C(n3410), .Y(n3394) );
  NAND3X1 U6645 ( .A(n3201), .B(n3208), .C(n3214), .Y(n3199) );
  NAND3X1 U6646 ( .A(n3162), .B(n3169), .C(n3175), .Y(n3160) );
  NAND3X1 U6647 ( .A(n3123), .B(n3130), .C(n3136), .Y(n3121) );
  NAND3X1 U6648 ( .A(n3079), .B(n3086), .C(n3093), .Y(n3077) );
  NAND3X1 U6649 ( .A(n2884), .B(n2891), .C(n2897), .Y(n2882) );
  NAND3X1 U6650 ( .A(n2845), .B(n2852), .C(n2858), .Y(n2843) );
  NAND3X1 U6651 ( .A(n2806), .B(n2813), .C(n2819), .Y(n2804) );
  NAND3X1 U6652 ( .A(n2762), .B(n2769), .C(n2776), .Y(n2760) );
  NAND3X1 U6653 ( .A(n2567), .B(n2574), .C(n2580), .Y(n2565) );
  NAND3X1 U6654 ( .A(n2528), .B(n2535), .C(n2541), .Y(n2526) );
  NAND3X1 U6655 ( .A(n2489), .B(n2496), .C(n2502), .Y(n2487) );
  NAND3X1 U6656 ( .A(n2445), .B(n2452), .C(n2459), .Y(n2443) );
  NAND3X1 U6657 ( .A(n2250), .B(n2257), .C(n2263), .Y(n2248) );
  NAND3X1 U6658 ( .A(n2211), .B(n2218), .C(n2224), .Y(n2209) );
  NAND3X1 U6659 ( .A(n2172), .B(n2179), .C(n2185), .Y(n2170) );
  NAND3X1 U6660 ( .A(n2128), .B(n2135), .C(n2142), .Y(n2126) );
  NAND3X1 U6661 ( .A(n2009), .B(n2014), .C(n2016), .Y(n2007) );
  NAND3X1 U6662 ( .A(n1970), .B(n1975), .C(n1977), .Y(n1968) );
  NAND3X1 U6663 ( .A(n1931), .B(n1936), .C(n1938), .Y(n1929) );
  NAND3X1 U6664 ( .A(n1892), .B(n1897), .C(n1899), .Y(n1890) );
  NAND3X1 U6665 ( .A(n1853), .B(n1858), .C(n1860), .Y(n1851) );
  NAND3X1 U6666 ( .A(n1809), .B(n1814), .C(n1816), .Y(n1807) );
  NAND3X1 U6667 ( .A(n1764), .B(n1769), .C(n1771), .Y(n1762) );
  NAND3X1 U6668 ( .A(n1720), .B(n1725), .C(n1727), .Y(n1718) );
  NAND3X1 U6669 ( .A(n1676), .B(n1681), .C(n1683), .Y(n1674) );
  NAND3X1 U6670 ( .A(n1632), .B(n1637), .C(n1639), .Y(n1630) );
  NAND3X1 U6671 ( .A(n1588), .B(n1593), .C(n1595), .Y(n1586) );
  NAND3X1 U6672 ( .A(n1544), .B(n1549), .C(n1551), .Y(n1542) );
  NAND3X1 U6673 ( .A(n1500), .B(n1505), .C(n1507), .Y(n1498) );
  AND3X2 U6674 ( .A(n1765), .B(n1771), .C(n5822), .Y(n1767) );
  AND3X2 U6675 ( .A(n1721), .B(n1727), .C(n5823), .Y(n1723) );
  AND3X2 U6676 ( .A(n1677), .B(n1683), .C(n5827), .Y(n1679) );
  AND3X2 U6677 ( .A(n1633), .B(n1639), .C(n5823), .Y(n1635) );
  AND3X2 U6678 ( .A(n1589), .B(n1595), .C(n5822), .Y(n1591) );
  AND3X2 U6679 ( .A(n1545), .B(n1551), .C(n5822), .Y(n1547) );
  AND3X2 U6680 ( .A(n1501), .B(n1507), .C(n5822), .Y(n1503) );
  AND3X2 U6681 ( .A(n1893), .B(n1899), .C(n5823), .Y(n1895) );
  AND3X2 U6682 ( .A(n1854), .B(n1860), .C(n5823), .Y(n1856) );
  OA22X2 U6683 ( .A0(n5851), .A1(n3950), .B0(n3957), .B1(n3952), .Y(n3933) );
  NOR2X1 U6684 ( .A(n3956), .B(n5799), .Y(n3957) );
  OA22X2 U6685 ( .A0(n5851), .A1(n3911), .B0(n3918), .B1(n3913), .Y(n3894) );
  NOR2X1 U6686 ( .A(n3917), .B(n5799), .Y(n3918) );
  OA22X2 U6687 ( .A0(n5853), .A1(n3872), .B0(n3879), .B1(n3874), .Y(n3855) );
  NOR2X1 U6688 ( .A(n3878), .B(n5799), .Y(n3879) );
  OA22X2 U6689 ( .A0(n5851), .A1(n3833), .B0(n3840), .B1(n3835), .Y(n3816) );
  NOR2X1 U6690 ( .A(n3839), .B(n5799), .Y(n3840) );
  OA22X2 U6691 ( .A0(n5851), .A1(n3794), .B0(n3801), .B1(n3796), .Y(n3777) );
  NOR2X1 U6692 ( .A(n3800), .B(n5799), .Y(n3801) );
  OA22X2 U6693 ( .A0(n5851), .A1(n3755), .B0(n3762), .B1(n3757), .Y(n3738) );
  NOR2X1 U6694 ( .A(n3761), .B(n5799), .Y(n3762) );
  OA22X2 U6695 ( .A0(n5851), .A1(n3711), .B0(n3718), .B1(n3713), .Y(n3694) );
  NOR2X1 U6696 ( .A(n3717), .B(n5799), .Y(n3718) );
  OA22X2 U6697 ( .A0(n5854), .A1(n3672), .B0(n3679), .B1(n3674), .Y(n3655) );
  NOR2X1 U6698 ( .A(n3678), .B(n5799), .Y(n3679) );
  OA22X2 U6699 ( .A0(n5854), .A1(n3633), .B0(n3640), .B1(n3635), .Y(n3616) );
  NOR2X1 U6700 ( .A(n3639), .B(n5800), .Y(n3640) );
  OA22X2 U6701 ( .A0(n5854), .A1(n3594), .B0(n3601), .B1(n3596), .Y(n3577) );
  NOR2X1 U6702 ( .A(n3600), .B(n5800), .Y(n3601) );
  OA22X2 U6703 ( .A0(n5854), .A1(n3555), .B0(n3562), .B1(n3557), .Y(n3538) );
  NOR2X1 U6704 ( .A(n3561), .B(n5800), .Y(n3562) );
  OA22X2 U6705 ( .A0(n5854), .A1(n3516), .B0(n3523), .B1(n3518), .Y(n3499) );
  NOR2X1 U6706 ( .A(n3522), .B(n5800), .Y(n3523) );
  OA22X2 U6707 ( .A0(n5854), .A1(n3477), .B0(n3484), .B1(n3479), .Y(n3460) );
  NOR2X1 U6708 ( .A(n3483), .B(n5800), .Y(n3484) );
  OA22X2 U6709 ( .A0(n5854), .A1(n3438), .B0(n3445), .B1(n3440), .Y(n3421) );
  NOR2X1 U6710 ( .A(n3444), .B(n5800), .Y(n3445) );
  OA22X2 U6711 ( .A0(n5854), .A1(n3394), .B0(n3401), .B1(n3396), .Y(n3377) );
  NOR2X1 U6712 ( .A(n3400), .B(n5800), .Y(n3401) );
  OA22X2 U6713 ( .A0(n5854), .A1(n3355), .B0(n3362), .B1(n3357), .Y(n3338) );
  NOR2X1 U6714 ( .A(n3361), .B(n5801), .Y(n3362) );
  OA22X2 U6715 ( .A0(n5854), .A1(n3316), .B0(n3323), .B1(n3318), .Y(n3299) );
  NOR2X1 U6716 ( .A(n3322), .B(n5801), .Y(n3323) );
  OA22X2 U6717 ( .A0(n5854), .A1(n3277), .B0(n3284), .B1(n3279), .Y(n3260) );
  NOR2X1 U6718 ( .A(n3283), .B(n5801), .Y(n3284) );
  OA22X2 U6719 ( .A0(n5854), .A1(n3238), .B0(n3245), .B1(n3240), .Y(n3221) );
  NOR2X1 U6720 ( .A(n3244), .B(n5801), .Y(n3245) );
  OA22X2 U6721 ( .A0(n5854), .A1(n3199), .B0(n3206), .B1(n3201), .Y(n3182) );
  NOR2X1 U6722 ( .A(n3205), .B(n5801), .Y(n3206) );
  OA22X2 U6723 ( .A0(n5854), .A1(n3160), .B0(n3167), .B1(n3162), .Y(n3143) );
  NOR2X1 U6724 ( .A(n3166), .B(n5801), .Y(n3167) );
  OA22X2 U6725 ( .A0(n5854), .A1(n3121), .B0(n3128), .B1(n3123), .Y(n3104) );
  NOR2X1 U6726 ( .A(n3127), .B(n5801), .Y(n3128) );
  OA22X2 U6727 ( .A0(n5854), .A1(n3077), .B0(n3084), .B1(n3079), .Y(n3060) );
  NOR2X1 U6728 ( .A(n3083), .B(n5801), .Y(n3084) );
  OA22X2 U6729 ( .A0(n5854), .A1(n3038), .B0(n3045), .B1(n3040), .Y(n3021) );
  NOR2X1 U6730 ( .A(n3044), .B(n5802), .Y(n3045) );
  OA22X2 U6731 ( .A0(n5854), .A1(n2999), .B0(n3006), .B1(n3001), .Y(n2982) );
  NOR2X1 U6732 ( .A(n3005), .B(n5802), .Y(n3006) );
  OA22X2 U6733 ( .A0(n5854), .A1(n2960), .B0(n2967), .B1(n2962), .Y(n2943) );
  NOR2X1 U6734 ( .A(n2966), .B(n5802), .Y(n2967) );
  OA22X2 U6735 ( .A0(n5853), .A1(n2921), .B0(n2928), .B1(n2923), .Y(n2904) );
  NOR2X1 U6736 ( .A(n2927), .B(n5802), .Y(n2928) );
  OA22X2 U6737 ( .A0(n5853), .A1(n2882), .B0(n2889), .B1(n2884), .Y(n2865) );
  NOR2X1 U6738 ( .A(n2888), .B(n5802), .Y(n2889) );
  OA22X2 U6739 ( .A0(n5853), .A1(n2843), .B0(n2850), .B1(n2845), .Y(n2826) );
  NOR2X1 U6740 ( .A(n2849), .B(n5802), .Y(n2850) );
  OA22X2 U6741 ( .A0(n5853), .A1(n2804), .B0(n2811), .B1(n2806), .Y(n2787) );
  NOR2X1 U6742 ( .A(n2810), .B(n5803), .Y(n2811) );
  OA22X2 U6743 ( .A0(n5853), .A1(n2760), .B0(n2767), .B1(n2762), .Y(n2743) );
  NOR2X1 U6744 ( .A(n2766), .B(n5803), .Y(n2767) );
  OA22X2 U6745 ( .A0(n5852), .A1(n2087), .B0(n2094), .B1(n2089), .Y(n2070) );
  NOR2X1 U6746 ( .A(n2093), .B(n5802), .Y(n2094) );
  OA22X2 U6747 ( .A0(n5852), .A1(n2048), .B0(n2055), .B1(n2050), .Y(n2031) );
  NOR2X1 U6748 ( .A(n2054), .B(n5802), .Y(n2055) );
  OA22X2 U6749 ( .A0(n5853), .A1(n2565), .B0(n2572), .B1(n2567), .Y(n2548) );
  NOR2X1 U6750 ( .A(n2571), .B(n5804), .Y(n2572) );
  OA22X2 U6751 ( .A0(n5853), .A1(n2526), .B0(n2533), .B1(n2528), .Y(n2509) );
  NOR2X1 U6752 ( .A(n2532), .B(n5804), .Y(n2533) );
  OA22X2 U6753 ( .A0(n5853), .A1(n2487), .B0(n2494), .B1(n2489), .Y(n2470) );
  NOR2X1 U6754 ( .A(n2493), .B(n5803), .Y(n2494) );
  OA22X2 U6755 ( .A0(n5853), .A1(n2443), .B0(n2450), .B1(n2445), .Y(n2426) );
  NOR2X1 U6756 ( .A(n2449), .B(n5804), .Y(n2450) );
  OA22X2 U6757 ( .A0(n5853), .A1(n2248), .B0(n2255), .B1(n2250), .Y(n2231) );
  NOR2X1 U6758 ( .A(n2254), .B(n5803), .Y(n2255) );
  OA22X2 U6759 ( .A0(n5853), .A1(n2209), .B0(n2216), .B1(n2211), .Y(n2192) );
  NOR2X1 U6760 ( .A(n2215), .B(n5803), .Y(n2216) );
  OA22X2 U6761 ( .A0(n5852), .A1(n2170), .B0(n2177), .B1(n2172), .Y(n2153) );
  NOR2X1 U6762 ( .A(n2176), .B(n5802), .Y(n2177) );
  OA22X2 U6763 ( .A0(n5852), .A1(n2126), .B0(n2133), .B1(n2128), .Y(n2109) );
  NOR2X1 U6764 ( .A(n2132), .B(n5802), .Y(n2133) );
  OAI222X4 U6765 ( .A0(n5798), .A1(n1023), .B0(n1036), .B1(n1025), .C0(n1033), 
        .C1(n5819), .Y(n984) );
  OA21XL U6766 ( .A0(n6573), .A1(n5849), .B0(n5828), .Y(n1036) );
  INVX3 U6767 ( .A(n2006), .Y(n6474) );
  OAI222XL U6768 ( .A0(n5813), .A1(n2007), .B0(n2008), .B1(n2009), .C0(n5819), 
        .C1(n2010), .Y(n2006) );
  OA21XL U6769 ( .A0(n6532), .A1(n5844), .B0(n5839), .Y(n2008) );
  INVX3 U6770 ( .A(n1967), .Y(n6476) );
  OAI222XL U6771 ( .A0(n5813), .A1(n1968), .B0(n1969), .B1(n1970), .C0(n5819), 
        .C1(n1971), .Y(n1967) );
  OA21XL U6772 ( .A0(n6540), .A1(n5844), .B0(n5839), .Y(n1969) );
  INVX3 U6773 ( .A(n1928), .Y(n6478) );
  OAI222XL U6774 ( .A0(n5813), .A1(n1929), .B0(n1930), .B1(n1931), .C0(n5821), 
        .C1(n1932), .Y(n1928) );
  OA21XL U6775 ( .A0(n6548), .A1(n5844), .B0(n5839), .Y(n1930) );
  INVX3 U6776 ( .A(n1889), .Y(n6480) );
  OAI222XL U6777 ( .A0(n5813), .A1(n1890), .B0(n1891), .B1(n1892), .C0(n5815), 
        .C1(n1893), .Y(n1889) );
  OA21XL U6778 ( .A0(n6556), .A1(n5844), .B0(n5841), .Y(n1891) );
  INVX3 U6779 ( .A(n1850), .Y(n6482) );
  OAI222XL U6780 ( .A0(n5813), .A1(n1851), .B0(n1852), .B1(n1853), .C0(n5816), 
        .C1(n1854), .Y(n1850) );
  OA21XL U6781 ( .A0(n6564), .A1(n5844), .B0(n5842), .Y(n1852) );
  INVX3 U6782 ( .A(n1806), .Y(n6484) );
  OAI222XL U6783 ( .A0(n5813), .A1(n1807), .B0(n1808), .B1(n1809), .C0(n5819), 
        .C1(n1810), .Y(n1806) );
  OA21XL U6784 ( .A0(n6572), .A1(n5850), .B0(n5828), .Y(n1808) );
  INVX3 U6785 ( .A(n3949), .Y(n6424) );
  OAI222XL U6786 ( .A0(n5808), .A1(n3950), .B0(n3951), .B1(n3952), .C0(n5821), 
        .C1(n3953), .Y(n3949) );
  OA21XL U6787 ( .A0(n6518), .A1(n5844), .B0(n5828), .Y(n3951) );
  INVX3 U6788 ( .A(n3910), .Y(n6425) );
  OAI222XL U6789 ( .A0(n5809), .A1(n3911), .B0(n3912), .B1(n3913), .C0(n5821), 
        .C1(n3914), .Y(n3910) );
  OA21XL U6790 ( .A0(n6526), .A1(n5844), .B0(n5837), .Y(n3912) );
  INVX3 U6791 ( .A(n3871), .Y(n6426) );
  OAI222XL U6792 ( .A0(n5813), .A1(n3872), .B0(n3873), .B1(n3874), .C0(n5821), 
        .C1(n3875), .Y(n3871) );
  OA21XL U6793 ( .A0(n6534), .A1(n5850), .B0(n5841), .Y(n3873) );
  INVX3 U6794 ( .A(n3832), .Y(n6427) );
  OAI222XL U6795 ( .A0(n5811), .A1(n3833), .B0(n3834), .B1(n3835), .C0(n5821), 
        .C1(n3836), .Y(n3832) );
  OA21XL U6796 ( .A0(n6542), .A1(n5849), .B0(n5828), .Y(n3834) );
  INVX3 U6797 ( .A(n3793), .Y(n6428) );
  OAI222XL U6798 ( .A0(n5813), .A1(n3794), .B0(n3795), .B1(n3796), .C0(n5821), 
        .C1(n3797), .Y(n3793) );
  OA21XL U6799 ( .A0(n6550), .A1(n5850), .B0(n5842), .Y(n3795) );
  INVX3 U6800 ( .A(n3754), .Y(n6429) );
  OAI222XL U6801 ( .A0(n5810), .A1(n3755), .B0(n3756), .B1(n3757), .C0(n5820), 
        .C1(n3758), .Y(n3754) );
  OA21XL U6802 ( .A0(n6558), .A1(n5850), .B0(n5840), .Y(n3756) );
  INVX3 U6803 ( .A(n3710), .Y(n6430) );
  OAI222XL U6804 ( .A0(n5812), .A1(n3711), .B0(n3712), .B1(n3713), .C0(n5821), 
        .C1(n3714), .Y(n3710) );
  OA21XL U6805 ( .A0(n6566), .A1(n5844), .B0(n5842), .Y(n3712) );
  INVX3 U6806 ( .A(n3671), .Y(n6431) );
  OAI222XL U6807 ( .A0(n5811), .A1(n3672), .B0(n3673), .B1(n3674), .C0(n5820), 
        .C1(n3675), .Y(n3671) );
  OA21XL U6808 ( .A0(n6511), .A1(n5849), .B0(n5842), .Y(n3673) );
  INVX3 U6809 ( .A(n3632), .Y(n6432) );
  OAI222XL U6810 ( .A0(n5811), .A1(n3633), .B0(n3634), .B1(n3635), .C0(n5820), 
        .C1(n3636), .Y(n3632) );
  OA21XL U6811 ( .A0(n6519), .A1(n5849), .B0(n5842), .Y(n3634) );
  INVX3 U6812 ( .A(n3593), .Y(n6433) );
  OAI222XL U6813 ( .A0(n5811), .A1(n3594), .B0(n3595), .B1(n3596), .C0(n5820), 
        .C1(n3597), .Y(n3593) );
  OA21XL U6814 ( .A0(n6527), .A1(n5849), .B0(n5842), .Y(n3595) );
  INVX3 U6815 ( .A(n3554), .Y(n6434) );
  OAI222XL U6816 ( .A0(n5811), .A1(n3555), .B0(n3556), .B1(n3557), .C0(n5819), 
        .C1(n3558), .Y(n3554) );
  OA21XL U6817 ( .A0(n6535), .A1(n5849), .B0(n5842), .Y(n3556) );
  INVX3 U6818 ( .A(n3515), .Y(n6435) );
  OAI222XL U6819 ( .A0(n5811), .A1(n3516), .B0(n3517), .B1(n3518), .C0(n5819), 
        .C1(n3519), .Y(n3515) );
  OA21XL U6820 ( .A0(n6543), .A1(n5844), .B0(n5842), .Y(n3517) );
  INVX3 U6821 ( .A(n3476), .Y(n6436) );
  OAI222XL U6822 ( .A0(n5811), .A1(n3477), .B0(n3478), .B1(n3479), .C0(n5820), 
        .C1(n3480), .Y(n3476) );
  OA21XL U6823 ( .A0(n6551), .A1(n5850), .B0(n5842), .Y(n3478) );
  INVX3 U6824 ( .A(n3437), .Y(n6437) );
  OAI222XL U6825 ( .A0(n5812), .A1(n3438), .B0(n3439), .B1(n3440), .C0(n5820), 
        .C1(n3441), .Y(n3437) );
  OA21XL U6826 ( .A0(n6559), .A1(n5849), .B0(n5830), .Y(n3439) );
  INVX3 U6827 ( .A(n3393), .Y(n6438) );
  OAI222XL U6828 ( .A0(n5811), .A1(n3394), .B0(n3395), .B1(n3396), .C0(n5819), 
        .C1(n3397), .Y(n3393) );
  OA21XL U6829 ( .A0(n6567), .A1(n5849), .B0(n5842), .Y(n3395) );
  INVX3 U6830 ( .A(n3354), .Y(n6439) );
  OAI222XL U6831 ( .A0(n5812), .A1(n3355), .B0(n3356), .B1(n3357), .C0(n5819), 
        .C1(n3358), .Y(n3354) );
  OA21XL U6832 ( .A0(n6512), .A1(n5850), .B0(n5839), .Y(n3356) );
  INVX3 U6833 ( .A(n3315), .Y(n6440) );
  OAI222XL U6834 ( .A0(n5813), .A1(n3316), .B0(n3317), .B1(n3318), .C0(n5819), 
        .C1(n3319), .Y(n3315) );
  OA21XL U6835 ( .A0(n6520), .A1(n5850), .B0(n5840), .Y(n3317) );
  INVX3 U6836 ( .A(n3276), .Y(n6441) );
  OAI222XL U6837 ( .A0(n5814), .A1(n3277), .B0(n3278), .B1(n3279), .C0(n5820), 
        .C1(n3280), .Y(n3276) );
  OA21XL U6838 ( .A0(n6528), .A1(n5850), .B0(n5837), .Y(n3278) );
  INVX3 U6839 ( .A(n3237), .Y(n6442) );
  OAI222XL U6840 ( .A0(n5812), .A1(n3238), .B0(n3239), .B1(n3240), .C0(n5819), 
        .C1(n3241), .Y(n3237) );
  OA21XL U6841 ( .A0(n6536), .A1(n5850), .B0(n5839), .Y(n3239) );
  INVX3 U6842 ( .A(n3198), .Y(n6443) );
  OAI222XL U6843 ( .A0(n5812), .A1(n3199), .B0(n3200), .B1(n3201), .C0(n5819), 
        .C1(n3202), .Y(n3198) );
  OA21XL U6844 ( .A0(n6544), .A1(n5850), .B0(n5841), .Y(n3200) );
  INVX3 U6845 ( .A(n3159), .Y(n6444) );
  OAI222XL U6846 ( .A0(n5812), .A1(n3160), .B0(n3161), .B1(n3162), .C0(n5819), 
        .C1(n3163), .Y(n3159) );
  OA21XL U6847 ( .A0(n6552), .A1(n5850), .B0(n5841), .Y(n3161) );
  INVX3 U6848 ( .A(n3120), .Y(n6445) );
  OAI222XL U6849 ( .A0(n5812), .A1(n3121), .B0(n3122), .B1(n3123), .C0(n5820), 
        .C1(n3124), .Y(n3120) );
  OA21XL U6850 ( .A0(n6560), .A1(n5850), .B0(n5841), .Y(n3122) );
  INVX3 U6851 ( .A(n3076), .Y(n6446) );
  OAI222XL U6852 ( .A0(n5812), .A1(n3077), .B0(n3078), .B1(n3079), .C0(n5819), 
        .C1(n3080), .Y(n3076) );
  OA21XL U6853 ( .A0(n6568), .A1(n5850), .B0(n5841), .Y(n3078) );
  INVX3 U6854 ( .A(n3037), .Y(n6447) );
  OAI222XL U6855 ( .A0(n5812), .A1(n3038), .B0(n3039), .B1(n3040), .C0(n5819), 
        .C1(n3041), .Y(n3037) );
  OA21XL U6856 ( .A0(n6513), .A1(n5844), .B0(n5841), .Y(n3039) );
  INVX3 U6857 ( .A(n2998), .Y(n6448) );
  OAI222XL U6858 ( .A0(n5812), .A1(n2999), .B0(n3000), .B1(n3001), .C0(n5820), 
        .C1(n3002), .Y(n2998) );
  OA21XL U6859 ( .A0(n6521), .A1(n5844), .B0(n5841), .Y(n3000) );
  INVX3 U6860 ( .A(n2959), .Y(n6449) );
  OAI222XL U6861 ( .A0(n5812), .A1(n2960), .B0(n2961), .B1(n2962), .C0(n5819), 
        .C1(n2963), .Y(n2959) );
  OA21XL U6862 ( .A0(n6529), .A1(n5844), .B0(n5841), .Y(n2961) );
  INVX3 U6863 ( .A(n2920), .Y(n6450) );
  OAI222XL U6864 ( .A0(n5813), .A1(n2921), .B0(n2922), .B1(n2923), .C0(n5819), 
        .C1(n2924), .Y(n2920) );
  OA21XL U6865 ( .A0(n6537), .A1(n5844), .B0(n5841), .Y(n2922) );
  INVX3 U6866 ( .A(n2881), .Y(n6451) );
  OAI222XL U6867 ( .A0(n5811), .A1(n2882), .B0(n2883), .B1(n2884), .C0(n5820), 
        .C1(n2885), .Y(n2881) );
  OA21XL U6868 ( .A0(n6545), .A1(n5844), .B0(n5841), .Y(n2883) );
  INVX3 U6869 ( .A(n2842), .Y(n6452) );
  OAI222XL U6870 ( .A0(n5812), .A1(n2843), .B0(n2844), .B1(n2845), .C0(n5820), 
        .C1(n2846), .Y(n2842) );
  OA21XL U6871 ( .A0(n6553), .A1(n5844), .B0(n5842), .Y(n2844) );
  INVX3 U6872 ( .A(n2803), .Y(n6453) );
  OAI222XL U6873 ( .A0(n5814), .A1(n2804), .B0(n2805), .B1(n2806), .C0(n5820), 
        .C1(n2807), .Y(n2803) );
  OA21XL U6874 ( .A0(n6561), .A1(n5844), .B0(n5840), .Y(n2805) );
  INVX3 U6875 ( .A(n2759), .Y(n6454) );
  OAI222XL U6876 ( .A0(n5811), .A1(n2760), .B0(n2761), .B1(n2762), .C0(n5820), 
        .C1(n2763), .Y(n2759) );
  OA21XL U6877 ( .A0(n6569), .A1(n5844), .B0(n5840), .Y(n2761) );
  INVX3 U6878 ( .A(n2086), .Y(n6471) );
  OAI222XL U6879 ( .A0(n5814), .A1(n2087), .B0(n2088), .B1(n2089), .C0(n5821), 
        .C1(n2090), .Y(n2086) );
  OA21XL U6880 ( .A0(n6516), .A1(n5849), .B0(n5839), .Y(n2088) );
  INVX3 U6881 ( .A(n2047), .Y(n6472) );
  OAI222XL U6882 ( .A0(n5811), .A1(n2048), .B0(n2049), .B1(n2050), .C0(n5819), 
        .C1(n2051), .Y(n2047) );
  OA21XL U6883 ( .A0(n6524), .A1(n5844), .B0(n5839), .Y(n2049) );
  INVX3 U6884 ( .A(n2564), .Y(n6459) );
  OAI222XL U6885 ( .A0(n5813), .A1(n2565), .B0(n2566), .B1(n2567), .C0(n5820), 
        .C1(n2568), .Y(n2564) );
  OA21XL U6886 ( .A0(n6546), .A1(n5849), .B0(n5840), .Y(n2566) );
  INVX3 U6887 ( .A(n2525), .Y(n6460) );
  OAI222XL U6888 ( .A0(n5814), .A1(n2526), .B0(n2527), .B1(n2528), .C0(n5821), 
        .C1(n2529), .Y(n2525) );
  OA21XL U6889 ( .A0(n6554), .A1(n5844), .B0(n5840), .Y(n2527) );
  INVX3 U6890 ( .A(n2486), .Y(n6461) );
  OAI222XL U6891 ( .A0(n5812), .A1(n2487), .B0(n2488), .B1(n2489), .C0(n5820), 
        .C1(n2490), .Y(n2486) );
  OA21XL U6892 ( .A0(n6562), .A1(n5849), .B0(n5840), .Y(n2488) );
  INVX3 U6893 ( .A(n2442), .Y(n6462) );
  OAI222XL U6894 ( .A0(n5814), .A1(n2443), .B0(n2444), .B1(n2445), .C0(n5821), 
        .C1(n2446), .Y(n2442) );
  OA21XL U6895 ( .A0(n6570), .A1(n5850), .B0(n5840), .Y(n2444) );
  INVX3 U6896 ( .A(n2247), .Y(n6467) );
  OAI222XL U6897 ( .A0(n5811), .A1(n2248), .B0(n2249), .B1(n2250), .C0(n5821), 
        .C1(n2251), .Y(n2247) );
  OA21XL U6898 ( .A0(n6547), .A1(n5850), .B0(n5828), .Y(n2249) );
  INVX3 U6899 ( .A(n2208), .Y(n6468) );
  OAI222XL U6900 ( .A0(n5813), .A1(n2209), .B0(n2210), .B1(n2211), .C0(n5821), 
        .C1(n2212), .Y(n2208) );
  OA21XL U6901 ( .A0(n6555), .A1(n5843), .B0(n5828), .Y(n2210) );
  INVX3 U6902 ( .A(n2169), .Y(n6469) );
  OAI222XL U6903 ( .A0(n5812), .A1(n2170), .B0(n2171), .B1(n2172), .C0(n5821), 
        .C1(n2173), .Y(n2169) );
  OA21XL U6904 ( .A0(n6563), .A1(n5843), .B0(n5828), .Y(n2171) );
  INVX3 U6905 ( .A(n2125), .Y(n6470) );
  OAI222XL U6906 ( .A0(n5814), .A1(n2126), .B0(n2127), .B1(n2128), .C0(n5821), 
        .C1(n2129), .Y(n2125) );
  OA21XL U6907 ( .A0(n6571), .A1(n5844), .B0(n5828), .Y(n2127) );
  AO22X2 U6908 ( .A0(n2091), .A1(n5765), .B0(n6516), .B1(n2095), .Y(n2068) );
  AO22X1 U6909 ( .A0(n2089), .A1(n5833), .B0(n2090), .B1(n5823), .Y(n2095) );
  AO22X2 U6910 ( .A0(n2052), .A1(n5765), .B0(n6524), .B1(n2056), .Y(n2029) );
  AO22X1 U6911 ( .A0(n2050), .A1(n5833), .B0(n2051), .B1(n5825), .Y(n2056) );
  CLKINVX1 U6912 ( .A(n4040), .Y(n6575) );
  CLKINVX1 U6913 ( .A(n3952), .Y(n6583) );
  CLKINVX1 U6914 ( .A(n3913), .Y(n6591) );
  CLKINVX1 U6915 ( .A(n3874), .Y(n6599) );
  CLKINVX1 U6916 ( .A(n3674), .Y(n6576) );
  CLKINVX1 U6917 ( .A(n3635), .Y(n6584) );
  CLKINVX1 U6918 ( .A(n3596), .Y(n6592) );
  CLKINVX1 U6919 ( .A(n3557), .Y(n6600) );
  CLKINVX1 U6920 ( .A(n3318), .Y(n6585) );
  CLKINVX1 U6921 ( .A(n3240), .Y(n6601) );
  CLKINVX1 U6922 ( .A(n3001), .Y(n6586) );
  CLKINVX1 U6923 ( .A(n2923), .Y(n6602) );
  CLKINVX1 U6924 ( .A(n2684), .Y(n6587) );
  CLKINVX1 U6925 ( .A(n2606), .Y(n6603) );
  CLKINVX1 U6926 ( .A(n2367), .Y(n6588) );
  CLKINVX1 U6927 ( .A(n2289), .Y(n6604) );
  CLKINVX1 U6928 ( .A(n2050), .Y(n6589) );
  CLKINVX1 U6929 ( .A(n3835), .Y(n6607) );
  CLKINVX1 U6930 ( .A(n3796), .Y(n6615) );
  CLKINVX1 U6931 ( .A(n3757), .Y(n6623) );
  CLKINVX1 U6932 ( .A(n3713), .Y(n6631) );
  CLKINVX1 U6933 ( .A(n3518), .Y(n6608) );
  CLKINVX1 U6934 ( .A(n3479), .Y(n6616) );
  CLKINVX1 U6935 ( .A(n3440), .Y(n6624) );
  CLKINVX1 U6936 ( .A(n3396), .Y(n6632) );
  BUFX4 U6937 ( .A(n5916), .Y(n5913) );
  BUFX4 U6938 ( .A(n5912), .Y(n5915) );
  BUFX4 U6939 ( .A(n5912), .Y(n5914) );
  AND2X2 U6940 ( .A(n1028), .B(n5807), .Y(n4827) );
  CLKINVX1 U6941 ( .A(n3357), .Y(n6577) );
  CLKINVX1 U6942 ( .A(n3279), .Y(n6593) );
  CLKINVX1 U6943 ( .A(n3040), .Y(n6578) );
  CLKINVX1 U6944 ( .A(n2962), .Y(n6594) );
  CLKINVX1 U6945 ( .A(n2723), .Y(n6579) );
  CLKINVX1 U6946 ( .A(n2645), .Y(n6595) );
  CLKINVX1 U6947 ( .A(n2406), .Y(n6580) );
  CLKINVX1 U6948 ( .A(n2328), .Y(n6596) );
  CLKINVX1 U6949 ( .A(n2089), .Y(n6581) );
  CLKINVX1 U6950 ( .A(n3201), .Y(n6609) );
  CLKINVX1 U6951 ( .A(n3162), .Y(n6617) );
  CLKINVX1 U6952 ( .A(n3123), .Y(n6625) );
  CLKINVX1 U6953 ( .A(n3079), .Y(n6633) );
  CLKINVX1 U6954 ( .A(n2884), .Y(n6610) );
  CLKINVX1 U6955 ( .A(n2845), .Y(n6618) );
  CLKINVX1 U6956 ( .A(n2806), .Y(n6626) );
  CLKINVX1 U6957 ( .A(n2762), .Y(n6634) );
  CLKINVX1 U6958 ( .A(n2567), .Y(n6611) );
  CLKINVX1 U6959 ( .A(n2528), .Y(n6619) );
  CLKINVX1 U6960 ( .A(n2489), .Y(n6627) );
  CLKINVX1 U6961 ( .A(n2445), .Y(n6635) );
  CLKINVX1 U6962 ( .A(n2250), .Y(n6612) );
  CLKINVX1 U6963 ( .A(n2211), .Y(n6620) );
  CLKINVX1 U6964 ( .A(n2172), .Y(n6628) );
  CLKINVX1 U6965 ( .A(n2128), .Y(n6636) );
  CLKINVX1 U6966 ( .A(n1025), .Y(n6638) );
  CLKINVX1 U6967 ( .A(n1764), .Y(n6582) );
  CLKINVX1 U6968 ( .A(n1720), .Y(n6590) );
  CLKINVX1 U6969 ( .A(n1676), .Y(n6598) );
  CLKINVX1 U6970 ( .A(n1632), .Y(n6606) );
  CLKINVX1 U6971 ( .A(n2009), .Y(n6597) );
  CLKINVX1 U6972 ( .A(n1970), .Y(n6605) );
  CLKINVX1 U6973 ( .A(n1931), .Y(n6613) );
  CLKINVX1 U6974 ( .A(n1892), .Y(n6621) );
  CLKINVX1 U6975 ( .A(n1853), .Y(n6629) );
  CLKINVX1 U6976 ( .A(n1809), .Y(n6637) );
  CLKINVX1 U6977 ( .A(n1588), .Y(n6614) );
  CLKINVX1 U6978 ( .A(n1544), .Y(n6622) );
  CLKINVX1 U6979 ( .A(n1500), .Y(n6630) );
  CLKBUFX3 U6980 ( .A(n5826), .Y(n5824) );
  CLKBUFX3 U6981 ( .A(n5826), .Y(n5825) );
  INVX3 U6982 ( .A(n5843), .Y(n5848) );
  NOR2X1 U6983 ( .A(n6646), .B(n6651), .Y(n974) );
  NAND2X1 U6984 ( .A(n5955), .B(n6651), .Y(n4083) );
  INVX3 U6985 ( .A(n3891), .Y(n6348) );
  INVX3 U6986 ( .A(n3813), .Y(n6350) );
  INVX3 U6987 ( .A(n3774), .Y(n6351) );
  INVX3 U6988 ( .A(n3613), .Y(n6355) );
  INVX3 U6989 ( .A(n3574), .Y(n6356) );
  INVX3 U6990 ( .A(n3535), .Y(n6357) );
  INVX3 U6991 ( .A(n3496), .Y(n6358) );
  INVX3 U6992 ( .A(n3457), .Y(n6359) );
  INVX3 U6993 ( .A(n3418), .Y(n6360) );
  INVX3 U6994 ( .A(n3374), .Y(n6361) );
  INVX3 U6995 ( .A(n3335), .Y(n6362) );
  INVX3 U6996 ( .A(n3296), .Y(n6363) );
  INVX3 U6997 ( .A(n3257), .Y(n6364) );
  INVX3 U6998 ( .A(n3218), .Y(n6365) );
  INVX3 U6999 ( .A(n3179), .Y(n6366) );
  INVX3 U7000 ( .A(n4674), .Y(n6367) );
  INVX3 U7001 ( .A(n3101), .Y(n6368) );
  INVX3 U7002 ( .A(n3057), .Y(n6369) );
  INVX3 U7003 ( .A(n3018), .Y(n6370) );
  INVX3 U7004 ( .A(n2979), .Y(n6371) );
  INVX3 U7005 ( .A(n4675), .Y(n6372) );
  INVX3 U7006 ( .A(n2901), .Y(n6373) );
  INVX3 U7007 ( .A(n2862), .Y(n6374) );
  INVX3 U7008 ( .A(n2823), .Y(n6375) );
  INVX3 U7009 ( .A(n2784), .Y(n6376) );
  INVX3 U7010 ( .A(n2740), .Y(n6377) );
  INVX3 U7011 ( .A(n2701), .Y(n6378) );
  INVX3 U7012 ( .A(n2662), .Y(n6379) );
  INVX3 U7013 ( .A(n2623), .Y(n6380) );
  INVX3 U7014 ( .A(n2584), .Y(n6381) );
  INVX3 U7015 ( .A(n2545), .Y(n6382) );
  INVX3 U7016 ( .A(n2506), .Y(n6383) );
  INVX3 U7017 ( .A(n2467), .Y(n6384) );
  INVX3 U7018 ( .A(n2423), .Y(n6385) );
  INVX3 U7019 ( .A(n2384), .Y(n6386) );
  INVX3 U7020 ( .A(n2345), .Y(n6387) );
  INVX3 U7021 ( .A(n2306), .Y(n6388) );
  INVX3 U7022 ( .A(n2267), .Y(n6389) );
  INVX3 U7023 ( .A(n2228), .Y(n6390) );
  INVX3 U7024 ( .A(n2189), .Y(n6391) );
  INVX3 U7025 ( .A(n2150), .Y(n6392) );
  INVX3 U7026 ( .A(n2106), .Y(n6393) );
  INVX3 U7027 ( .A(n2067), .Y(n6394) );
  INVX3 U7028 ( .A(n2028), .Y(n6395) );
  INVX3 U7029 ( .A(n1949), .Y(n6397) );
  INVX3 U7030 ( .A(n1699), .Y(n6402) );
  INVX3 U7031 ( .A(n1655), .Y(n6403) );
  INVX3 U7032 ( .A(n1611), .Y(n6404) );
  INVX3 U7033 ( .A(n1567), .Y(n6405) );
  INVX3 U7034 ( .A(n1523), .Y(n6406) );
  INVX3 U7035 ( .A(n1479), .Y(n6407) );
  CLKBUFX3 U7036 ( .A(n4669), .Y(n5761) );
  CLKBUFX3 U7037 ( .A(n4669), .Y(n5762) );
  CLKBUFX3 U7038 ( .A(n4669), .Y(n5763) );
  INVX3 U7039 ( .A(n5756), .Y(n5754) );
  CLKBUFX3 U7040 ( .A(n4814), .Y(n5756) );
  INVX3 U7041 ( .A(n4814), .Y(n5753) );
  INVX3 U7042 ( .A(n5757), .Y(n5752) );
  CLKBUFX3 U7043 ( .A(n4814), .Y(n5757) );
  INVX3 U7044 ( .A(n5796), .Y(n5794) );
  INVX3 U7045 ( .A(n5870), .Y(n5869) );
  INVX3 U7046 ( .A(n5882), .Y(n5879) );
  CLKINVX1 U7047 ( .A(n5660), .Y(n6227) );
  CLKINVX1 U7048 ( .A(n5665), .Y(n6194) );
  CLKBUFX3 U7049 ( .A(n5959), .Y(n5456) );
  CLKBUFX3 U7050 ( .A(n5924), .Y(n5923) );
  CLKINVX1 U7051 ( .A(n5660), .Y(n6258) );
  CLKINVX1 U7052 ( .A(n5657), .Y(n6036) );
  CLKINVX1 U7053 ( .A(n5657), .Y(n6066) );
  CLKINVX1 U7054 ( .A(n5657), .Y(n6003) );
  CLKBUFX3 U7055 ( .A(n5969), .Y(n5065) );
  NAND2X2 U7056 ( .A(n5667), .B(n3961), .Y(n3722) );
  INVX6 U7057 ( .A(n5937), .Y(n5935) );
  CLKBUFX3 U7058 ( .A(n5939), .Y(n5937) );
  INVX6 U7059 ( .A(n5942), .Y(n5941) );
  CLKBUFX3 U7060 ( .A(n5943), .Y(n5942) );
  CLKBUFX3 U7061 ( .A(n5269), .Y(n5268) );
  CLKBUFX3 U7062 ( .A(n5933), .Y(n5931) );
  CLKINVX1 U7063 ( .A(N3358), .Y(n6131) );
  CLKINVX1 U7064 ( .A(N3358), .Y(n6098) );
  CLKINVX1 U7065 ( .A(n4667), .Y(n6132) );
  CLKINVX1 U7066 ( .A(n4667), .Y(n6099) );
  CLKINVX1 U7067 ( .A(n4667), .Y(n6162) );
  CLKINVX1 U7068 ( .A(N3353), .Y(n6133) );
  CLKINVX1 U7069 ( .A(N3353), .Y(n6100) );
  CLKINVX1 U7070 ( .A(N3353), .Y(n6163) );
  CLKINVX1 U7071 ( .A(N3360), .Y(n6260) );
  CLKINVX1 U7072 ( .A(N3360), .Y(n6195) );
  CLKINVX1 U7073 ( .A(N3360), .Y(n6228) );
  CLKBUFX3 U7074 ( .A(n5933), .Y(n5932) );
  INVX6 U7075 ( .A(n5919), .Y(n5917) );
  CLKBUFX3 U7076 ( .A(n4668), .Y(n5949) );
  INVX3 U7077 ( .A(n4884), .Y(n5858) );
  INVX3 U7078 ( .A(n4886), .Y(n5875) );
  INVX3 U7079 ( .A(n4884), .Y(n5855) );
  INVX3 U7080 ( .A(n4884), .Y(n5856) );
  INVX3 U7081 ( .A(n4884), .Y(n5857) );
  INVX3 U7082 ( .A(n4885), .Y(n5863) );
  INVX3 U7083 ( .A(n4885), .Y(n5864) );
  INVX3 U7084 ( .A(n4885), .Y(n5865) );
  INVX3 U7085 ( .A(n4886), .Y(n5872) );
  INVX3 U7086 ( .A(n4886), .Y(n5873) );
  INVX3 U7087 ( .A(n4886), .Y(n5874) );
  INVX3 U7088 ( .A(n4887), .Y(n5883) );
  INVX3 U7089 ( .A(n4887), .Y(n5884) );
  INVX3 U7090 ( .A(n4887), .Y(n5885) );
  INVX3 U7091 ( .A(n4888), .Y(n5893) );
  INVX3 U7092 ( .A(n4888), .Y(n5894) );
  INVX3 U7093 ( .A(n4888), .Y(n5895) );
  INVX3 U7094 ( .A(n4889), .Y(n5903) );
  INVX3 U7095 ( .A(n4889), .Y(n5904) );
  INVX3 U7096 ( .A(n4889), .Y(n5905) );
  INVX3 U7097 ( .A(n4890), .Y(n5909) );
  INVX3 U7098 ( .A(n4890), .Y(n5910) );
  INVX3 U7099 ( .A(n4890), .Y(n5911) );
  INVX3 U7100 ( .A(n4891), .Y(n5906) );
  INVX3 U7101 ( .A(n4891), .Y(n5907) );
  INVX3 U7102 ( .A(n4891), .Y(n5908) );
  CLKBUFX3 U7103 ( .A(n6508), .Y(n5746) );
  CLKINVX1 U7104 ( .A(n5664), .Y(n6507) );
  CLKBUFX3 U7105 ( .A(n6505), .Y(n5734) );
  CLKINVX1 U7106 ( .A(n5661), .Y(n6505) );
  CLKBUFX3 U7107 ( .A(n6506), .Y(n5737) );
  CLKBUFX3 U7108 ( .A(n6503), .Y(n5727) );
  CLKINVX1 U7109 ( .A(N3360), .Y(n6503) );
  CLKBUFX3 U7110 ( .A(n6504), .Y(n5731) );
  CLKBUFX3 U7111 ( .A(n4893), .Y(n5270) );
  CLKINVX1 U7112 ( .A(n5658), .Y(n6101) );
  CLKINVX1 U7113 ( .A(n5658), .Y(n6165) );
  CLKINVX1 U7114 ( .A(n5651), .Y(n6007) );
  CLKINVX1 U7115 ( .A(n5651), .Y(n6070) );
  NOR2BX1 U7116 ( .AN(n4061), .B(n1476), .Y(n966) );
  INVX6 U7117 ( .A(n5927), .Y(n5925) );
  AND2X2 U7118 ( .A(n1441), .B(n1430), .Y(n4061) );
  NOR3BX2 U7119 ( .AN(n4666), .B(n5955), .C(N3327), .Y(n3097) );
  NOR3BX2 U7120 ( .AN(n4666), .B(n5270), .C(N3327), .Y(n2780) );
  NOR3BX2 U7121 ( .AN(n4666), .B(n6639), .C(n5955), .Y(n3731) );
  NOR3BX2 U7122 ( .AN(n4666), .B(n6639), .C(n5270), .Y(n3414) );
  NAND2X2 U7123 ( .A(n3732), .B(n1785), .Y(n4040) );
  NAND2X2 U7124 ( .A(n3732), .B(n1740), .Y(n3952) );
  NAND2X2 U7125 ( .A(n3732), .B(n1696), .Y(n3913) );
  NAND2X2 U7126 ( .A(n3732), .B(n1652), .Y(n3874) );
  NAND2X2 U7127 ( .A(n3732), .B(n1608), .Y(n3835) );
  NAND2X2 U7128 ( .A(n3732), .B(n1564), .Y(n3796) );
  NAND2X2 U7129 ( .A(n3732), .B(n1520), .Y(n3757) );
  NAND2X2 U7130 ( .A(n3732), .B(n1066), .Y(n3713) );
  NAND2X2 U7131 ( .A(n3415), .B(n1785), .Y(n3674) );
  NAND2X2 U7132 ( .A(n3415), .B(n1740), .Y(n3635) );
  NAND2X2 U7133 ( .A(n3415), .B(n1696), .Y(n3596) );
  NAND2X2 U7134 ( .A(n3415), .B(n1652), .Y(n3557) );
  NAND2X2 U7135 ( .A(n3415), .B(n1608), .Y(n3518) );
  NAND2X2 U7136 ( .A(n3415), .B(n1564), .Y(n3479) );
  NAND2X2 U7137 ( .A(n3415), .B(n1520), .Y(n3440) );
  NAND2X2 U7138 ( .A(n3415), .B(n1066), .Y(n3396) );
  NAND2X2 U7139 ( .A(n3098), .B(n1740), .Y(n3318) );
  NAND2X2 U7140 ( .A(n3098), .B(n1652), .Y(n3240) );
  NAND2X2 U7141 ( .A(n2781), .B(n1740), .Y(n3001) );
  NAND2X2 U7142 ( .A(n2781), .B(n1652), .Y(n2923) );
  NAND2X2 U7143 ( .A(n2464), .B(n1740), .Y(n2684) );
  NAND2X2 U7144 ( .A(n2464), .B(n1652), .Y(n2606) );
  NAND2X2 U7145 ( .A(n2147), .B(n1740), .Y(n2367) );
  NAND2X2 U7146 ( .A(n2147), .B(n1652), .Y(n2289) );
  NAND2X2 U7147 ( .A(n1829), .B(n1740), .Y(n2050) );
  INVX6 U7148 ( .A(n5938), .Y(n5934) );
  CLKBUFX3 U7149 ( .A(n5939), .Y(n5938) );
  INVX6 U7150 ( .A(n5943), .Y(n5940) );
  CLKBUFX3 U7151 ( .A(n5827), .Y(n5822) );
  CLKBUFX3 U7152 ( .A(n5797), .Y(n5807) );
  CLKBUFX3 U7153 ( .A(n5829), .Y(n5835) );
  CLKBUFX3 U7154 ( .A(n5912), .Y(n5916) );
  CLKBUFX3 U7155 ( .A(n6417), .Y(n5678) );
  NAND2X2 U7156 ( .A(n3098), .B(n1785), .Y(n3357) );
  NAND2X2 U7157 ( .A(n3098), .B(n1696), .Y(n3279) );
  NAND2X2 U7158 ( .A(n3098), .B(n1608), .Y(n3201) );
  NAND2X2 U7159 ( .A(n3098), .B(n1564), .Y(n3162) );
  NAND2X2 U7160 ( .A(n3098), .B(n1520), .Y(n3123) );
  NAND2X2 U7161 ( .A(n3098), .B(n1066), .Y(n3079) );
  NAND2X2 U7162 ( .A(n2781), .B(n1785), .Y(n3040) );
  NAND2X2 U7163 ( .A(n2781), .B(n1696), .Y(n2962) );
  NAND2X2 U7164 ( .A(n2781), .B(n1608), .Y(n2884) );
  NAND2X2 U7165 ( .A(n2781), .B(n1564), .Y(n2845) );
  NAND2X2 U7166 ( .A(n2781), .B(n1520), .Y(n2806) );
  NAND2X2 U7167 ( .A(n2781), .B(n1066), .Y(n2762) );
  NAND2X2 U7168 ( .A(n2464), .B(n1785), .Y(n2723) );
  NAND2X2 U7169 ( .A(n2464), .B(n1696), .Y(n2645) );
  NAND2X2 U7170 ( .A(n2147), .B(n1785), .Y(n2406) );
  NAND2X2 U7171 ( .A(n2147), .B(n1696), .Y(n2328) );
  NAND2X2 U7172 ( .A(n1829), .B(n1785), .Y(n2089) );
  NAND2X2 U7173 ( .A(n2464), .B(n1608), .Y(n2567) );
  NAND2X2 U7174 ( .A(n2464), .B(n1564), .Y(n2528) );
  NAND2X2 U7175 ( .A(n2464), .B(n1520), .Y(n2489) );
  NAND2X2 U7176 ( .A(n2464), .B(n1066), .Y(n2445) );
  NAND2X2 U7177 ( .A(n2147), .B(n1608), .Y(n2250) );
  NAND2X2 U7178 ( .A(n2147), .B(n1564), .Y(n2211) );
  NAND2X2 U7179 ( .A(n2147), .B(n1520), .Y(n2172) );
  NAND2X2 U7180 ( .A(n2147), .B(n1066), .Y(n2128) );
  CLKBUFX3 U7181 ( .A(n5827), .Y(n5823) );
  CLKBUFX3 U7182 ( .A(n5829), .Y(n5836) );
  CLKBUFX3 U7183 ( .A(n5829), .Y(n5837) );
  CLKBUFX3 U7184 ( .A(n5830), .Y(n5842) );
  CLKBUFX3 U7185 ( .A(n5830), .Y(n5841) );
  CLKBUFX3 U7186 ( .A(n5830), .Y(n5840) );
  CLKBUFX3 U7187 ( .A(n5830), .Y(n5839) );
  CLKBUFX3 U7188 ( .A(n5844), .Y(n5850) );
  CLKBUFX3 U7189 ( .A(n5843), .Y(n5849) );
  CLKBUFX3 U7190 ( .A(n5797), .Y(n5808) );
  CLKBUFX3 U7191 ( .A(n5808), .Y(n5810) );
  CLKBUFX3 U7192 ( .A(n5797), .Y(n5809) );
  CLKINVX1 U7193 ( .A(N3359), .Y(n6502) );
  CLKINVX1 U7194 ( .A(N3357), .Y(n6501) );
  CLKINVX1 U7195 ( .A(n5659), .Y(n6500) );
  AOI221XL U7196 ( .A0(n5270), .A1(n6651), .B0(n6646), .B1(n5955), .C0(n6645), 
        .Y(n4084) );
  CLKINVX1 U7197 ( .A(n4087), .Y(n6645) );
  CLKINVX1 U7198 ( .A(n4088), .Y(n6651) );
  CLKINVX1 U7199 ( .A(n4081), .Y(n6646) );
  CLKBUFX3 U7200 ( .A(n5798), .Y(n5811) );
  CLKBUFX3 U7201 ( .A(n5798), .Y(n5812) );
  CLKBUFX3 U7202 ( .A(n5798), .Y(n5813) );
  CLKBUFX3 U7203 ( .A(n5798), .Y(n5814) );
  CLKBUFX3 U7204 ( .A(n5837), .Y(n5838) );
  NAND2X2 U7205 ( .A(n5951), .B(n3496), .Y(n3495) );
  NAND2X2 U7206 ( .A(n5951), .B(n3457), .Y(n3456) );
  NAND2X2 U7207 ( .A(n5951), .B(n3418), .Y(n3417) );
  NAND2X2 U7208 ( .A(cur_state), .B(n3374), .Y(n3373) );
  NAND2X2 U7209 ( .A(n5951), .B(n3335), .Y(n3334) );
  NAND2X2 U7210 ( .A(cur_state), .B(n3296), .Y(n3295) );
  NAND2X2 U7211 ( .A(n5951), .B(n3257), .Y(n3256) );
  NAND2X2 U7212 ( .A(cur_state), .B(n3218), .Y(n3217) );
  NAND2X2 U7213 ( .A(n5951), .B(n3179), .Y(n3178) );
  NAND2X2 U7214 ( .A(n5951), .B(n3101), .Y(n3100) );
  NAND2X2 U7215 ( .A(cur_state), .B(n3057), .Y(n3056) );
  NAND2X2 U7216 ( .A(n5951), .B(n3018), .Y(n3017) );
  NAND2X2 U7217 ( .A(cur_state), .B(n2979), .Y(n2978) );
  NAND2X2 U7218 ( .A(n5951), .B(n2901), .Y(n2900) );
  NAND2X2 U7219 ( .A(cur_state), .B(n2862), .Y(n2861) );
  NAND2X2 U7220 ( .A(n5951), .B(n2823), .Y(n2822) );
  NAND2X2 U7221 ( .A(n5951), .B(n2784), .Y(n2783) );
  NAND2X2 U7222 ( .A(cur_state), .B(n2740), .Y(n2739) );
  NAND2X2 U7223 ( .A(n5951), .B(n2701), .Y(n2700) );
  NAND2X2 U7224 ( .A(cur_state), .B(n2623), .Y(n2622) );
  NAND2X2 U7225 ( .A(n5951), .B(n2584), .Y(n2583) );
  NAND2X2 U7226 ( .A(cur_state), .B(n2545), .Y(n2544) );
  NAND2X2 U7227 ( .A(cur_state), .B(n2506), .Y(n2505) );
  NAND2X2 U7228 ( .A(n5953), .B(n2467), .Y(n2466) );
  NAND2X2 U7229 ( .A(n5953), .B(n2423), .Y(n2422) );
  NAND2X2 U7230 ( .A(n5953), .B(n2384), .Y(n2383) );
  NAND2X2 U7231 ( .A(n5953), .B(n2345), .Y(n2344) );
  NAND2X2 U7232 ( .A(n5953), .B(n2306), .Y(n2305) );
  NAND2X2 U7233 ( .A(n5953), .B(n2267), .Y(n2266) );
  NAND2X2 U7234 ( .A(n5953), .B(n2228), .Y(n2227) );
  NAND2X2 U7235 ( .A(n5953), .B(n2189), .Y(n2188) );
  NAND2X2 U7236 ( .A(n5953), .B(n2150), .Y(n2149) );
  NAND2X2 U7237 ( .A(n5953), .B(n2106), .Y(n2105) );
  NAND2X2 U7238 ( .A(cur_state), .B(n2067), .Y(n2066) );
  NAND2X2 U7239 ( .A(n5951), .B(n2028), .Y(n2027) );
  NAND2X2 U7240 ( .A(n5951), .B(n1949), .Y(n1948) );
  NAND2X2 U7241 ( .A(cur_state), .B(n1699), .Y(n1698) );
  NAND2X2 U7242 ( .A(n5951), .B(n1655), .Y(n1654) );
  NAND2X2 U7243 ( .A(cur_state), .B(n1611), .Y(n1610) );
  OA22X4 U7244 ( .A0(n1980), .A1(n4627), .B0(n1643), .B1(n1820), .Y(n4830) );
  OA22X4 U7245 ( .A0(n1941), .A1(n4627), .B0(n1599), .B1(n1820), .Y(n4831) );
  OA22X4 U7246 ( .A0(n1902), .A1(n4627), .B0(n1555), .B1(n1820), .Y(n4832) );
  AOI221XL U7247 ( .A0(n3982), .A1(n5658), .B0(n3983), .B1(n5948), .C0(n3984), 
        .Y(n3974) );
  AOI221XL U7248 ( .A0(N3353), .A1(n3982), .B0(n5944), .B1(n3983), .C0(n3995), 
        .Y(n3992) );
  MX4X1 U7249 ( .A(n5291), .B(n5289), .C(n5290), .D(n5288), .S0(n4800), .S1(
        n5959), .Y(n5292) );
  MX4X1 U7250 ( .A(n5281), .B(n5279), .C(n5280), .D(n5278), .S0(n4800), .S1(
        n5959), .Y(n5282) );
  BUFX12 U7251 ( .A(N3365), .Y(n5664) );
  MX4X1 U7252 ( .A(n5331), .B(n5329), .C(n5330), .D(n5328), .S0(n4800), .S1(
        n5959), .Y(n5332) );
  MX4X1 U7253 ( .A(n5321), .B(n5319), .C(n5320), .D(n5318), .S0(n4800), .S1(
        n5959), .Y(n5322) );
  INVX3 U7254 ( .A(n5795), .Y(n5793) );
  CLKBUFX3 U7255 ( .A(n5796), .Y(n5795) );
  INVX3 U7256 ( .A(n5871), .Y(n5866) );
  INVX3 U7257 ( .A(n5871), .Y(n5867) );
  INVX3 U7258 ( .A(n5870), .Y(n5868) );
  CLKBUFX3 U7259 ( .A(n5871), .Y(n5870) );
  INVX3 U7260 ( .A(n5882), .Y(n5876) );
  INVX3 U7261 ( .A(n5881), .Y(n5877) );
  CLKBUFX3 U7262 ( .A(n5882), .Y(n5881) );
  INVX3 U7263 ( .A(n5880), .Y(n5878) );
  CLKBUFX3 U7264 ( .A(n5882), .Y(n5880) );
  INVX3 U7265 ( .A(n5892), .Y(n5886) );
  INVX3 U7266 ( .A(n5892), .Y(n5887) );
  INVX3 U7267 ( .A(n5891), .Y(n5888) );
  CLKBUFX3 U7268 ( .A(n5892), .Y(n5891) );
  INVX3 U7269 ( .A(n5902), .Y(n5896) );
  INVX3 U7270 ( .A(n5901), .Y(n5897) );
  CLKBUFX3 U7271 ( .A(n5902), .Y(n5901) );
  INVX3 U7272 ( .A(n5900), .Y(n5898) );
  CLKBUFX3 U7273 ( .A(n5902), .Y(n5900) );
  OA22X4 U7274 ( .A0(n2731), .A1(n4627), .B0(n1775), .B1(n2454), .Y(n4837) );
  OA22X4 U7275 ( .A0(n2692), .A1(n4627), .B0(n1731), .B1(n2454), .Y(n4838) );
  OA22X4 U7276 ( .A0(n2653), .A1(n4627), .B0(n1687), .B1(n2454), .Y(n4839) );
  OA22X4 U7277 ( .A0(n2614), .A1(n4627), .B0(n1643), .B1(n2454), .Y(n4840) );
  OA22X4 U7278 ( .A0(n2575), .A1(n4627), .B0(n1599), .B1(n2454), .Y(n4841) );
  OA22X4 U7279 ( .A0(n2536), .A1(n4627), .B0(n1555), .B1(n2454), .Y(n4842) );
  OA22X4 U7280 ( .A0(n2497), .A1(n4627), .B0(n1511), .B1(n2454), .Y(n4843) );
  OA22X4 U7281 ( .A0(n2453), .A1(n4627), .B0(n1042), .B1(n2454), .Y(n4844) );
  OA22X4 U7282 ( .A0(n2414), .A1(n4627), .B0(n1775), .B1(n2137), .Y(n4845) );
  OA22X4 U7283 ( .A0(n2375), .A1(n4627), .B0(n1731), .B1(n2137), .Y(n4846) );
  OA22X4 U7284 ( .A0(n2336), .A1(n4627), .B0(n1687), .B1(n2137), .Y(n4847) );
  OA22X4 U7285 ( .A0(n2297), .A1(n4627), .B0(n1643), .B1(n2137), .Y(n4848) );
  OA22X4 U7286 ( .A0(n2258), .A1(n4627), .B0(n1599), .B1(n2137), .Y(n4849) );
  OA22X4 U7287 ( .A0(n2219), .A1(n4627), .B0(n1555), .B1(n2137), .Y(n4850) );
  OA22X4 U7288 ( .A0(n2180), .A1(n4627), .B0(n1511), .B1(n2137), .Y(n4851) );
  OA22X4 U7289 ( .A0(n2136), .A1(n4627), .B0(n1042), .B1(n2137), .Y(n4852) );
  OA22X4 U7290 ( .A0(n2097), .A1(n4627), .B0(n1775), .B1(n1820), .Y(n4853) );
  OA22X4 U7291 ( .A0(n2058), .A1(n4627), .B0(n1731), .B1(n1820), .Y(n4854) );
  OA22X4 U7292 ( .A0(n3682), .A1(n4627), .B0(n1775), .B1(n3405), .Y(n4855) );
  OA22X4 U7293 ( .A0(n3643), .A1(n4627), .B0(n1731), .B1(n3405), .Y(n4856) );
  OA22X4 U7294 ( .A0(n3604), .A1(n4627), .B0(n1687), .B1(n3405), .Y(n4857) );
  OA22X4 U7295 ( .A0(n3565), .A1(n4627), .B0(n1643), .B1(n3405), .Y(n4858) );
  OA22X4 U7296 ( .A0(n3526), .A1(n4627), .B0(n1599), .B1(n3405), .Y(n4859) );
  OA22X4 U7297 ( .A0(n3487), .A1(n4627), .B0(n1555), .B1(n3405), .Y(n4860) );
  OA22X4 U7298 ( .A0(n3448), .A1(n4627), .B0(n1511), .B1(n3405), .Y(n4861) );
  OA22X4 U7299 ( .A0(n3404), .A1(n4627), .B0(n1042), .B1(n3405), .Y(n4862) );
  OA22X4 U7300 ( .A0(n3365), .A1(n4627), .B0(n1775), .B1(n3088), .Y(n4863) );
  OA22X4 U7301 ( .A0(n3326), .A1(n4627), .B0(n1731), .B1(n3088), .Y(n4864) );
  OA22X4 U7302 ( .A0(n3287), .A1(n4627), .B0(n1687), .B1(n3088), .Y(n4865) );
  OA22X4 U7303 ( .A0(n3248), .A1(n4627), .B0(n1643), .B1(n3088), .Y(n4866) );
  OA22X4 U7304 ( .A0(n3209), .A1(n4627), .B0(n1599), .B1(n3088), .Y(n4867) );
  OA22X4 U7305 ( .A0(n3131), .A1(n4627), .B0(n1511), .B1(n3088), .Y(n4868) );
  OA22X4 U7306 ( .A0(n3087), .A1(n4627), .B0(n1042), .B1(n3088), .Y(n4869) );
  OA22X4 U7307 ( .A0(n3048), .A1(n4627), .B0(n1775), .B1(n2771), .Y(n4870) );
  OA22X4 U7308 ( .A0(n3009), .A1(n4627), .B0(n1731), .B1(n2771), .Y(n4871) );
  OA22X4 U7309 ( .A0(n2931), .A1(n4627), .B0(n1643), .B1(n2771), .Y(n4872) );
  OA22X4 U7310 ( .A0(n2892), .A1(n4627), .B0(n1599), .B1(n2771), .Y(n4873) );
  OA22X4 U7311 ( .A0(n2853), .A1(n4627), .B0(n1555), .B1(n2771), .Y(n4874) );
  OA22X4 U7312 ( .A0(n2814), .A1(n4627), .B0(n1511), .B1(n2771), .Y(n4875) );
  OA22X4 U7313 ( .A0(n2770), .A1(n4627), .B0(n1042), .B1(n2771), .Y(n4876) );
  OA22X4 U7314 ( .A0(n3960), .A1(n4627), .B0(n1731), .B1(n3722), .Y(n4878) );
  OA22X4 U7315 ( .A0(n3921), .A1(n4627), .B0(n1687), .B1(n3722), .Y(n4879) );
  OA22X4 U7316 ( .A0(n3882), .A1(n4627), .B0(n1643), .B1(n3722), .Y(n4880) );
  OA22X4 U7317 ( .A0(n3843), .A1(n4627), .B0(n1599), .B1(n3722), .Y(n4881) );
  OA22X4 U7318 ( .A0(n3804), .A1(n4627), .B0(n1555), .B1(n3722), .Y(n4882) );
  MX4X1 U7319 ( .A(n5141), .B(n5139), .C(n5140), .D(n5138), .S0(n5272), .S1(
        n5267), .Y(n5142) );
  MX4X1 U7320 ( .A(n5131), .B(n5129), .C(n5130), .D(n5128), .S0(n5272), .S1(
        n5267), .Y(n5132) );
  MX4X1 U7321 ( .A(n5091), .B(n5089), .C(n5090), .D(n5088), .S0(n5272), .S1(
        n5647), .Y(n5092) );
  MX4X1 U7322 ( .A(n5086), .B(n5084), .C(n5085), .D(n5083), .S0(n5272), .S1(
        n5647), .Y(n5087) );
  MX4X1 U7323 ( .A(n4898), .B(n4896), .C(n4897), .D(n4895), .S0(n5067), .S1(
        n5065), .Y(n4899) );
  MX4X1 U7324 ( .A(n4908), .B(n4906), .C(n4907), .D(n4905), .S0(n5067), .S1(
        n5065), .Y(n4909) );
  MX4X1 U7325 ( .A(n4983), .B(n4981), .C(n4982), .D(n4980), .S0(n5068), .S1(
        n5969), .Y(n4984) );
  CLKBUFX3 U7326 ( .A(N3348), .Y(n5655) );
  MX4X1 U7327 ( .A(n4974), .B(n4964), .C(n4969), .D(n4959), .S0(N3322), .S1(
        N3321), .Y(N3348) );
  MX4X1 U7328 ( .A(n5522), .B(n5520), .C(n5521), .D(n5519), .S0(n5648), .S1(
        n5269), .Y(n5523) );
  NAND2X1 U7329 ( .A(n5952), .B(n6642), .Y(n1040) );
  CLKINVX1 U7330 ( .A(N3339), .Y(n4892) );
  MX4X1 U7331 ( .A(n5121), .B(n5119), .C(n5120), .D(n5118), .S0(n5272), .S1(
        n5267), .Y(n5122) );
  MX4X1 U7332 ( .A(n5111), .B(n5109), .C(n5110), .D(n5108), .S0(n5272), .S1(
        n5268), .Y(n5112) );
  MX4X1 U7333 ( .A(n5202), .B(n5192), .C(n5197), .D(n5187), .S0(n4666), .S1(
        N3327), .Y(N3354) );
  MX4X1 U7334 ( .A(n5201), .B(n5199), .C(n5200), .D(n5198), .S0(n5271), .S1(
        n5268), .Y(n5202) );
  MX4X1 U7335 ( .A(n5181), .B(n5179), .C(n5180), .D(n5178), .S0(n5271), .S1(
        n5268), .Y(n5182) );
  MX4X1 U7336 ( .A(n5171), .B(n5169), .C(n5170), .D(n5168), .S0(n5271), .S1(
        n5267), .Y(n5172) );
  MX4X1 U7337 ( .A(n5161), .B(n5159), .C(n5160), .D(n5158), .S0(n5271), .S1(
        n5267), .Y(n5162) );
  MX4X1 U7338 ( .A(n5151), .B(n5149), .C(n5150), .D(n5148), .S0(n5271), .S1(
        n5267), .Y(n5152) );
  INVX3 U7339 ( .A(reset), .Y(n6642) );
  CLKBUFX3 U7340 ( .A(n1776), .Y(n5667) );
  NOR2X1 U7341 ( .A(n5954), .B(reset), .Y(n1776) );
  MX4X1 U7342 ( .A(n5603), .B(n5593), .C(n5598), .D(n5588), .S0(n5672), .S1(
        n5674), .Y(n5463) );
  MX4X1 U7343 ( .A(n5602), .B(n5600), .C(n5601), .D(n5599), .S0(n5649), .S1(
        n5963), .Y(n5603) );
  MX4X1 U7344 ( .A(n5543), .B(n5533), .C(n5538), .D(n5528), .S0(n5672), .S1(
        n5674), .Y(n5460) );
  MX4X1 U7345 ( .A(n5583), .B(n5573), .C(n5578), .D(n5568), .S0(n5672), .S1(
        n5674), .Y(n5462) );
  OAI21X2 U7346 ( .A0(n5953), .A1(n971), .B0(n6642), .Y(n967) );
  NOR2BX1 U7347 ( .AN(n967), .B(reset), .Y(n4093) );
  NOR2X2 U7348 ( .A(n5671), .B(reset), .Y(n1068) );
  AOI2BB1X1 U7349 ( .A0N(reset), .A1N(n4087), .B0(n6641), .Y(n4086) );
  AO21X1 U7350 ( .A0(n4088), .A1(n4082), .B0(n6641), .Y(n4085) );
  NOR2X2 U7351 ( .A(n4000), .B(n4627), .Y(N16287) );
  OAI2BB2XL U7352 ( .B0(n4094), .B1(n6658), .A0N(N3454), .A1N(n4095), .Y(n4621) );
  OAI2BB2XL U7353 ( .B0(n4094), .B1(n6657), .A0N(N3453), .A1N(n4095), .Y(n4622) );
  OAI2BB2XL U7354 ( .B0(n4094), .B1(n6656), .A0N(N3452), .A1N(n4095), .Y(n4623) );
  OAI2BB2XL U7355 ( .B0(n4094), .B1(n6655), .A0N(N3451), .A1N(n4095), .Y(n4624) );
  OAI2BB2XL U7356 ( .B0(n6664), .B1(n967), .A0N(N3384), .A1N(n4093), .Y(n4615)
         );
  OAI2BB2XL U7357 ( .B0(n6662), .B1(n967), .A0N(N3382), .A1N(n4093), .Y(n4617)
         );
  OAI2BB2XL U7358 ( .B0(n6663), .B1(n967), .A0N(N3383), .A1N(n4093), .Y(n4616)
         );
  OAI2BB2XL U7359 ( .B0(n6661), .B1(n967), .A0N(N3381), .A1N(n4093), .Y(n4618)
         );
  OAI22XL U7360 ( .A0(n6641), .A1(n4089), .B0(n4819), .B1(n4080), .Y(n4613) );
  AOI211X1 U7361 ( .A0(n6650), .A1(N3339), .B0(n4090), .C0(reset), .Y(n4089)
         );
  CLKINVX1 U7362 ( .A(n4083), .Y(n6650) );
  AOI31X1 U7363 ( .A0(n4088), .A1(n6666), .A2(n4084), .B0(n4819), .Y(n4090) );
  CLKINVX1 U7364 ( .A(n4080), .Y(n6641) );
  OAI22XL U7365 ( .A0(n5964), .A1(n4064), .B0(reset), .B1(n4065), .Y(n4609) );
  OAI31XL U7366 ( .A0(n4068), .A1(n5253), .A2(n6665), .B0(n6652), .Y(n4066) );
  CLKINVX1 U7367 ( .A(n4069), .Y(n6652) );
  OAI22XL U7368 ( .A0(n5078), .A1(n4064), .B0(reset), .B1(n4070), .Y(n4610) );
  AOI21X1 U7369 ( .A0(n5634), .A1(n4071), .B0(n4072), .Y(n4070) );
  AOI211X1 U7370 ( .A0(n6665), .A1(n4073), .B0(n5250), .C0(n6640), .Y(n4072)
         );
  CLKINVX1 U7371 ( .A(n4064), .Y(n6640) );
  AND2X1 U7372 ( .A(n4094), .B(n6642), .Y(n4095) );
  OAI21XL U7373 ( .A0(n4077), .A1(n6666), .B0(n4078), .Y(n4611) );
  NAND4X1 U7374 ( .A(n4079), .B(n4080), .C(n6642), .D(n6666), .Y(n4078) );
  AOI2BB1X1 U7375 ( .A0N(n4084), .A1N(reset), .B0(n6641), .Y(n4077) );
  OAI31XL U7376 ( .A0(n4081), .A1(n5955), .A2(n4082), .B0(n4083), .Y(n4079) );
  CLKBUFX3 U7377 ( .A(N3352), .Y(n5658) );
  MX4X1 U7378 ( .A(n5242), .B(n5232), .C(n5237), .D(n5227), .S0(n4666), .S1(
        N3327), .Y(N3352) );
  MX4X1 U7379 ( .A(n5241), .B(n5239), .C(n5240), .D(n5238), .S0(n5270), .S1(
        n5268), .Y(n5242) );
  MX4X1 U7380 ( .A(n5231), .B(n5229), .C(n5230), .D(n5228), .S0(n5270), .S1(
        n5268), .Y(n5232) );
  NOR3X4 U7381 ( .A(n6655), .B(n6654), .C(n6656), .Y(n1430) );
  NOR3X4 U7382 ( .A(n6658), .B(n6657), .C(n6653), .Y(n1441) );
  NAND2X2 U7383 ( .A(n1475), .B(n1435), .Y(n1172) );
  NAND2X2 U7384 ( .A(n1470), .B(n1435), .Y(n1160) );
  NAND2X2 U7385 ( .A(n1446), .B(n1435), .Y(n1104) );
  NAND2X2 U7386 ( .A(n1428), .B(n1435), .Y(n1085) );
  NAND2X2 U7387 ( .A(n1475), .B(n1429), .Y(n1166) );
  NAND2X2 U7388 ( .A(n1470), .B(n1429), .Y(n1154) );
  NAND2X2 U7389 ( .A(n1446), .B(n1429), .Y(n1106) );
  NAND2X2 U7390 ( .A(n1428), .B(n1429), .Y(n1079) );
  NAND2X2 U7391 ( .A(n1451), .B(n1429), .Y(n1114) );
  NAND2X2 U7392 ( .A(n1446), .B(n1430), .Y(n1105) );
  NAND2X2 U7393 ( .A(n1428), .B(n1430), .Y(n1078) );
  NAND2X2 U7394 ( .A(n1470), .B(n1430), .Y(n1153) );
  NAND2X2 U7395 ( .A(n1475), .B(n1430), .Y(n1165) );
  NAND2X2 U7396 ( .A(n1435), .B(n1441), .Y(n1093) );
  NAND2X2 U7397 ( .A(n1429), .B(n1441), .Y(n1096) );
  NAND4X1 U7398 ( .A(n1452), .B(n1453), .C(n1454), .D(n1455), .Y(n1420) );
  NOR4X1 U7399 ( .A(n1466), .B(n1467), .C(n1468), .D(n1469), .Y(n1453) );
  NOR4X1 U7400 ( .A(n1461), .B(n1462), .C(n1463), .D(n1464), .Y(n1454) );
  NOR4X1 U7401 ( .A(n1471), .B(n1472), .C(n1473), .D(n1474), .Y(n1452) );
  NAND4X1 U7402 ( .A(n1399), .B(n1400), .C(n1401), .D(n1402), .Y(n1379) );
  NOR4X1 U7403 ( .A(n1411), .B(n1412), .C(n1413), .D(n1414), .Y(n1400) );
  NOR4X1 U7404 ( .A(n1407), .B(n1408), .C(n1409), .D(n1410), .Y(n1401) );
  NOR4X1 U7405 ( .A(n1415), .B(n1416), .C(n1417), .D(n1418), .Y(n1399) );
  NAND4X1 U7406 ( .A(n1358), .B(n1359), .C(n1360), .D(n1361), .Y(n1338) );
  NOR4X1 U7407 ( .A(n1370), .B(n1371), .C(n1372), .D(n1373), .Y(n1359) );
  NOR4X1 U7408 ( .A(n1366), .B(n1367), .C(n1368), .D(n1369), .Y(n1360) );
  NOR4X1 U7409 ( .A(n1374), .B(n1375), .C(n1376), .D(n1377), .Y(n1358) );
  NAND4X1 U7410 ( .A(n1317), .B(n1318), .C(n1319), .D(n1320), .Y(n1297) );
  NOR4X1 U7411 ( .A(n1329), .B(n1330), .C(n1331), .D(n1332), .Y(n1318) );
  NOR4X1 U7412 ( .A(n1325), .B(n1326), .C(n1327), .D(n1328), .Y(n1319) );
  NOR4X1 U7413 ( .A(n1333), .B(n1334), .C(n1335), .D(n1336), .Y(n1317) );
  NAND4X1 U7414 ( .A(n1276), .B(n1277), .C(n1278), .D(n1279), .Y(n1256) );
  NOR4X1 U7415 ( .A(n1288), .B(n1289), .C(n1290), .D(n1291), .Y(n1277) );
  NOR4X1 U7416 ( .A(n1284), .B(n1285), .C(n1286), .D(n1287), .Y(n1278) );
  NOR4X1 U7417 ( .A(n1292), .B(n1293), .C(n1294), .D(n1295), .Y(n1276) );
  NAND4X1 U7418 ( .A(n1235), .B(n1236), .C(n1237), .D(n1238), .Y(n1215) );
  NOR4X1 U7419 ( .A(n1247), .B(n1248), .C(n1249), .D(n1250), .Y(n1236) );
  NOR4X1 U7420 ( .A(n1243), .B(n1244), .C(n1245), .D(n1246), .Y(n1237) );
  NOR4X1 U7421 ( .A(n1251), .B(n1252), .C(n1253), .D(n1254), .Y(n1235) );
  NAND4X1 U7422 ( .A(n1121), .B(n1122), .C(n1123), .D(n1124), .Y(n1070) );
  NOR4X1 U7423 ( .A(n1149), .B(n1150), .C(n1151), .D(n1152), .Y(n1122) );
  NOR4X1 U7424 ( .A(n1137), .B(n1138), .C(n1139), .D(n1140), .Y(n1123) );
  NOR4X1 U7425 ( .A(n1161), .B(n1162), .C(n1163), .D(n1164), .Y(n1121) );
  NAND4X1 U7426 ( .A(n1194), .B(n1195), .C(n1196), .D(n1197), .Y(n1174) );
  NOR4X1 U7427 ( .A(n1206), .B(n1207), .C(n1208), .D(n1209), .Y(n1195) );
  NOR4X1 U7428 ( .A(n1202), .B(n1203), .C(n1204), .D(n1205), .Y(n1196) );
  NOR4X1 U7429 ( .A(n1210), .B(n1211), .C(n1212), .D(n1213), .Y(n1194) );
  NAND2X2 U7430 ( .A(n1451), .B(n1435), .Y(n1120) );
  NAND2X2 U7431 ( .A(n1451), .B(n1430), .Y(n1113) );
  NOR2BX1 U7432 ( .AN(n3961), .B(n1775), .Y(n971) );
  INVX3 U7433 ( .A(N3339), .Y(n6666) );
  NOR3X1 U7434 ( .A(n6664), .B(n6663), .C(n6659), .Y(n3961) );
  CLKBUFX3 U7435 ( .A(n1035), .Y(n5797) );
  CLKBUFX3 U7436 ( .A(n1031), .Y(n5829) );
  CLKBUFX3 U7437 ( .A(n1028), .Y(n5843) );
  NOR4X1 U7438 ( .A(n5764), .B(n5831), .C(n5822), .D(n6644), .Y(n976) );
  CLKINVX1 U7439 ( .A(n4000), .Y(n6644) );
  CLKBUFX3 U7440 ( .A(n1034), .Y(n5815) );
  NOR3X4 U7441 ( .A(n5270), .B(n5672), .C(n6666), .Y(n2464) );
  NOR3X4 U7442 ( .A(n5955), .B(n5672), .C(n6666), .Y(n2147) );
  NOR3X4 U7443 ( .A(n5966), .B(n5963), .C(n5964), .Y(n1608) );
  NOR3X4 U7444 ( .A(n5252), .B(n5963), .C(n5964), .Y(n1564) );
  NOR3X4 U7445 ( .A(n4749), .B(n5963), .C(n5966), .Y(n1520) );
  NOR3X4 U7446 ( .A(n4749), .B(n5963), .C(n5634), .Y(n1066) );
  CLKINVX1 U7447 ( .A(n3975), .Y(n6649) );
  CLKBUFX3 U7448 ( .A(n4748), .Y(n5964) );
  CLKBUFX3 U7449 ( .A(n1031), .Y(n5830) );
  CLKBUFX3 U7450 ( .A(n1031), .Y(n5828) );
  CLKBUFX3 U7451 ( .A(n1028), .Y(n5844) );
  CLKINVX1 U7452 ( .A(n4071), .Y(n6648) );
  AOI32X1 U7453 ( .A0(n5673), .A1(n6651), .A2(N3339), .B0(n4082), .B1(n6646), 
        .Y(n4087) );
  NAND2X1 U7454 ( .A(n4060), .B(n4057), .Y(n1476) );
  NAND2X1 U7455 ( .A(n4058), .B(n4059), .Y(n4068) );
  NAND2X1 U7456 ( .A(n4058), .B(n4060), .Y(n4088) );
  NOR2X1 U7457 ( .A(n5673), .B(N3339), .Y(n4082) );
  NAND2X1 U7458 ( .A(n4059), .B(n4057), .Y(n4081) );
  AND2X2 U7459 ( .A(n4068), .B(n4073), .Y(n975) );
  CLKBUFX3 U7460 ( .A(n1035), .Y(n5798) );
  CLKINVX1 U7461 ( .A(n4074), .Y(n6665) );
  OAI222XL U7462 ( .A0(n3933), .A1(n5724), .B0(n3934), .B1(n5701), .C0(n6424), 
        .C1(n5750), .Y(n3948) );
  OAI222XL U7463 ( .A0(n3894), .A1(n5724), .B0(n3895), .B1(n5699), .C0(n6425), 
        .C1(n5749), .Y(n3909) );
  OAI222XL U7464 ( .A0(n3855), .A1(n5724), .B0(n3856), .B1(n5698), .C0(n6426), 
        .C1(n5749), .Y(n3870) );
  OAI222XL U7465 ( .A0(n3816), .A1(n5724), .B0(n3817), .B1(n5698), .C0(n6427), 
        .C1(n5749), .Y(n3831) );
  OAI222XL U7466 ( .A0(n3777), .A1(n5724), .B0(n3778), .B1(n5698), .C0(n6428), 
        .C1(n5749), .Y(n3792) );
  OAI222XL U7467 ( .A0(n3738), .A1(n5724), .B0(n3739), .B1(n5701), .C0(n6429), 
        .C1(n5751), .Y(n3753) );
  OAI222XL U7468 ( .A0(n3694), .A1(n5724), .B0(n3695), .B1(n5701), .C0(n6430), 
        .C1(n5751), .Y(n3709) );
  OAI222XL U7469 ( .A0(n3655), .A1(n5724), .B0(n3656), .B1(n5698), .C0(n6431), 
        .C1(n5749), .Y(n3670) );
  OAI222XL U7470 ( .A0(n3616), .A1(n5724), .B0(n3617), .B1(n5698), .C0(n6432), 
        .C1(n6509), .Y(n3631) );
  OAI222XL U7471 ( .A0(n3577), .A1(n5724), .B0(n3578), .B1(n5698), .C0(n6433), 
        .C1(n6509), .Y(n3592) );
  OAI222XL U7472 ( .A0(n3538), .A1(n5724), .B0(n3539), .B1(n5698), .C0(n6434), 
        .C1(n5749), .Y(n3553) );
  OAI222XL U7473 ( .A0(n3499), .A1(n5725), .B0(n3500), .B1(n5701), .C0(n6435), 
        .C1(n5751), .Y(n3514) );
  OAI222XL U7474 ( .A0(n3460), .A1(n5725), .B0(n3461), .B1(n5700), .C0(n6436), 
        .C1(n5749), .Y(n3475) );
  OAI222XL U7475 ( .A0(n3421), .A1(n5725), .B0(n3422), .B1(n5700), .C0(n6437), 
        .C1(n5749), .Y(n3436) );
  OAI222XL U7476 ( .A0(n3377), .A1(n5725), .B0(n3378), .B1(n5700), .C0(n6438), 
        .C1(n5749), .Y(n3392) );
  OAI222XL U7477 ( .A0(n3338), .A1(n5725), .B0(n3339), .B1(n5700), .C0(n6439), 
        .C1(n5749), .Y(n3353) );
  OAI222XL U7478 ( .A0(n3299), .A1(n5725), .B0(n3300), .B1(n5701), .C0(n6440), 
        .C1(n5751), .Y(n3314) );
  OAI222XL U7479 ( .A0(n3260), .A1(n5725), .B0(n3261), .B1(n5701), .C0(n6441), 
        .C1(n5751), .Y(n3275) );
  OAI222XL U7480 ( .A0(n3221), .A1(n5725), .B0(n3222), .B1(n5701), .C0(n6442), 
        .C1(n5751), .Y(n3236) );
  OAI222XL U7481 ( .A0(n3182), .A1(n5725), .B0(n3183), .B1(n5701), .C0(n6443), 
        .C1(n5751), .Y(n3197) );
  OAI222XL U7482 ( .A0(n3143), .A1(n5725), .B0(n3144), .B1(n5701), .C0(n6444), 
        .C1(n5751), .Y(n3158) );
  OAI222XL U7483 ( .A0(n3104), .A1(n5725), .B0(n3105), .B1(n5701), .C0(n6445), 
        .C1(n5751), .Y(n3119) );
  OAI222XL U7484 ( .A0(n3060), .A1(n5725), .B0(n3061), .B1(n5701), .C0(n6446), 
        .C1(n5751), .Y(n3075) );
  OAI222XL U7485 ( .A0(n3021), .A1(n5726), .B0(n3022), .B1(n5701), .C0(n6447), 
        .C1(n5751), .Y(n3036) );
  OAI222XL U7486 ( .A0(n2982), .A1(n5726), .B0(n2983), .B1(n5701), .C0(n6448), 
        .C1(n5751), .Y(n2997) );
  OAI222XL U7487 ( .A0(n2943), .A1(n5726), .B0(n2944), .B1(n5701), .C0(n6449), 
        .C1(n5751), .Y(n2958) );
  OAI222XL U7488 ( .A0(n2904), .A1(n5726), .B0(n2905), .B1(n5701), .C0(n6450), 
        .C1(n5751), .Y(n2919) );
  OAI222XL U7489 ( .A0(n2865), .A1(n5726), .B0(n2866), .B1(n5701), .C0(n6451), 
        .C1(n5751), .Y(n2880) );
  OAI222XL U7490 ( .A0(n2826), .A1(n5726), .B0(n2827), .B1(n5701), .C0(n6452), 
        .C1(n5751), .Y(n2841) );
  OAI222XL U7491 ( .A0(n6376), .A1(n5856), .B0(n2801), .B1(n2783), .C0(n469), 
        .C1(n2784), .Y(n4367) );
  AOI211X1 U7492 ( .A0(n5917), .A1(n2785), .B0(n2802), .C0(n5792), .Y(n2801)
         );
  OAI222XL U7493 ( .A0(n2787), .A1(n5726), .B0(n2788), .B1(n5701), .C0(n6453), 
        .C1(n5751), .Y(n2802) );
  OAI222XL U7494 ( .A0(n6377), .A1(n5856), .B0(n2757), .B1(n2739), .C0(n461), 
        .C1(n2740), .Y(n4359) );
  AOI211X1 U7495 ( .A0(N3375), .A1(n2741), .B0(n2758), .C0(n5792), .Y(n2757)
         );
  OAI222XL U7496 ( .A0(n2743), .A1(n5726), .B0(n2744), .B1(n5701), .C0(n6454), 
        .C1(n5751), .Y(n2758) );
  OAI222XL U7497 ( .A0(n6378), .A1(n5856), .B0(n2718), .B1(n2700), .C0(n453), 
        .C1(n2701), .Y(n4351) );
  AOI211X1 U7498 ( .A0(n5917), .A1(n2702), .B0(n2719), .C0(n5792), .Y(n2718)
         );
  OAI222XL U7499 ( .A0(n2704), .A1(n5726), .B0(n2705), .B1(n5701), .C0(n6455), 
        .C1(n5751), .Y(n2719) );
  OAI222XL U7500 ( .A0(n6379), .A1(n5856), .B0(n2679), .B1(n2661), .C0(n445), 
        .C1(n2662), .Y(n4343) );
  AOI211X1 U7501 ( .A0(N3375), .A1(n2663), .B0(n2680), .C0(n5792), .Y(n2679)
         );
  OAI222XL U7502 ( .A0(n2665), .A1(n5726), .B0(n2666), .B1(n5700), .C0(n6456), 
        .C1(n5751), .Y(n2680) );
  OAI222XL U7503 ( .A0(n6380), .A1(n5856), .B0(n2640), .B1(n2622), .C0(n437), 
        .C1(n2623), .Y(n4335) );
  AOI211X1 U7504 ( .A0(n5917), .A1(n2624), .B0(n2641), .C0(n5792), .Y(n2640)
         );
  OAI222XL U7505 ( .A0(n2626), .A1(n5726), .B0(n2627), .B1(n5700), .C0(n6457), 
        .C1(n5749), .Y(n2641) );
  OAI222XL U7506 ( .A0(n6381), .A1(n5856), .B0(n2601), .B1(n2583), .C0(n429), 
        .C1(n2584), .Y(n4327) );
  AOI211X1 U7507 ( .A0(N3375), .A1(n2585), .B0(n2602), .C0(n5792), .Y(n2601)
         );
  OAI222XL U7508 ( .A0(n2587), .A1(n5726), .B0(n2588), .B1(n5700), .C0(n6458), 
        .C1(n5749), .Y(n2602) );
  OAI222XL U7509 ( .A0(n2548), .A1(n5726), .B0(n2549), .B1(n5700), .C0(n6459), 
        .C1(n5749), .Y(n2563) );
  OAI222XL U7510 ( .A0(n6383), .A1(n5857), .B0(n2523), .B1(n2505), .C0(n413), 
        .C1(n2506), .Y(n4311) );
  AOI211X1 U7511 ( .A0(n5917), .A1(n2507), .B0(n2524), .C0(n5792), .Y(n2523)
         );
  OAI222XL U7512 ( .A0(n2509), .A1(n5726), .B0(n2510), .B1(n5700), .C0(n6460), 
        .C1(n5749), .Y(n2524) );
  OAI222XL U7513 ( .A0(n6384), .A1(n5857), .B0(n2484), .B1(n2466), .C0(n405), 
        .C1(n2467), .Y(n4303) );
  AOI211X1 U7514 ( .A0(N3375), .A1(n2468), .B0(n2485), .C0(n5792), .Y(n2484)
         );
  OAI222XL U7515 ( .A0(n2470), .A1(n5726), .B0(n2471), .B1(n5700), .C0(n6461), 
        .C1(n5750), .Y(n2485) );
  OAI222XL U7516 ( .A0(n6385), .A1(n5857), .B0(n2440), .B1(n2422), .C0(n397), 
        .C1(n2423), .Y(n4295) );
  AOI211X1 U7517 ( .A0(N3375), .A1(n2424), .B0(n2441), .C0(n5793), .Y(n2440)
         );
  OAI222XL U7518 ( .A0(n2426), .A1(n5725), .B0(n2427), .B1(n5700), .C0(n6462), 
        .C1(n5750), .Y(n2441) );
  OAI222XL U7519 ( .A0(n6386), .A1(n5857), .B0(n2401), .B1(n2383), .C0(n389), 
        .C1(n2384), .Y(n4287) );
  AOI211X1 U7520 ( .A0(n5917), .A1(n2385), .B0(n2402), .C0(n5793), .Y(n2401)
         );
  OAI222XL U7521 ( .A0(n2387), .A1(n5725), .B0(n2388), .B1(n5700), .C0(n6463), 
        .C1(n5749), .Y(n2402) );
  OAI222XL U7522 ( .A0(n6387), .A1(n5857), .B0(n2362), .B1(n2344), .C0(n381), 
        .C1(n2345), .Y(n4279) );
  AOI211X1 U7523 ( .A0(N3375), .A1(n2346), .B0(n2363), .C0(n5793), .Y(n2362)
         );
  OAI222XL U7524 ( .A0(n2348), .A1(n5724), .B0(n2349), .B1(n5700), .C0(n6464), 
        .C1(n5750), .Y(n2363) );
  OAI222XL U7525 ( .A0(n6388), .A1(n5857), .B0(n2323), .B1(n2305), .C0(n373), 
        .C1(n2306), .Y(n4271) );
  AOI211X1 U7526 ( .A0(n5917), .A1(n2307), .B0(n2324), .C0(n5793), .Y(n2323)
         );
  OAI222XL U7527 ( .A0(n2309), .A1(n5726), .B0(n2310), .B1(n5700), .C0(n6465), 
        .C1(n5749), .Y(n2324) );
  OAI222XL U7528 ( .A0(n6389), .A1(n5857), .B0(n2284), .B1(n2266), .C0(n365), 
        .C1(n2267), .Y(n4263) );
  AOI211X1 U7529 ( .A0(N3375), .A1(n2268), .B0(n2285), .C0(n5793), .Y(n2284)
         );
  OAI222XL U7530 ( .A0(n2270), .A1(n6502), .B0(n2271), .B1(n5700), .C0(n6466), 
        .C1(n5750), .Y(n2285) );
  OAI222XL U7531 ( .A0(n6390), .A1(n5857), .B0(n2245), .B1(n2227), .C0(n357), 
        .C1(n2228), .Y(n4255) );
  AOI211X1 U7532 ( .A0(N3375), .A1(n2229), .B0(n2246), .C0(n5793), .Y(n2245)
         );
  OAI222XL U7533 ( .A0(n2231), .A1(n4824), .B0(n2232), .B1(n5700), .C0(n6467), 
        .C1(n6509), .Y(n2246) );
  OAI222XL U7534 ( .A0(n6391), .A1(n5857), .B0(n2206), .B1(n2188), .C0(n349), 
        .C1(n2189), .Y(n4247) );
  AOI211X1 U7535 ( .A0(n5917), .A1(n2190), .B0(n2207), .C0(n5793), .Y(n2206)
         );
  OAI222XL U7536 ( .A0(n2192), .A1(n5725), .B0(n2193), .B1(n5700), .C0(n6468), 
        .C1(n5749), .Y(n2207) );
  OAI222XL U7537 ( .A0(n6392), .A1(n5857), .B0(n2167), .B1(n2149), .C0(n341), 
        .C1(n2150), .Y(n4239) );
  AOI211X1 U7538 ( .A0(N3375), .A1(n2151), .B0(n2168), .C0(n5793), .Y(n2167)
         );
  OAI222XL U7539 ( .A0(n2153), .A1(n6502), .B0(n2154), .B1(n5700), .C0(n6469), 
        .C1(n6509), .Y(n2168) );
  OAI222XL U7540 ( .A0(n6393), .A1(n5857), .B0(n2123), .B1(n2105), .C0(n333), 
        .C1(n2106), .Y(n4231) );
  AOI211X1 U7541 ( .A0(n5917), .A1(n2107), .B0(n2124), .C0(n5793), .Y(n2123)
         );
  OAI222XL U7542 ( .A0(n2109), .A1(n5726), .B0(n2110), .B1(n5700), .C0(n6470), 
        .C1(n5749), .Y(n2124) );
  OAI222XL U7543 ( .A0(n6394), .A1(n5858), .B0(n2084), .B1(n2066), .C0(n325), 
        .C1(n2067), .Y(n4223) );
  AOI211X1 U7544 ( .A0(N3375), .A1(n2068), .B0(n2085), .C0(n5793), .Y(n2084)
         );
  OAI222XL U7545 ( .A0(n2070), .A1(n5725), .B0(n2071), .B1(n5700), .C0(n6471), 
        .C1(n5749), .Y(n2085) );
  OAI222XL U7546 ( .A0(n6395), .A1(n5858), .B0(n2045), .B1(n2027), .C0(n317), 
        .C1(n2028), .Y(n4215) );
  AOI211X1 U7547 ( .A0(n5917), .A1(n2029), .B0(n2046), .C0(n5793), .Y(n2045)
         );
  OAI222XL U7548 ( .A0(n2031), .A1(n5725), .B0(n2032), .B1(n5699), .C0(n6472), 
        .C1(n5749), .Y(n2046) );
  OAI222XL U7549 ( .A0(n6396), .A1(n5858), .B0(n2004), .B1(n1987), .C0(n309), 
        .C1(n1988), .Y(n4207) );
  AOI211X1 U7550 ( .A0(N3375), .A1(n6473), .B0(n2005), .C0(n5793), .Y(n2004)
         );
  OAI222XL U7551 ( .A0(n1990), .A1(n5726), .B0(n1991), .B1(n5699), .C0(n6474), 
        .C1(n5750), .Y(n2005) );
  OAI222XL U7552 ( .A0(n6397), .A1(n5858), .B0(n1965), .B1(n1948), .C0(n301), 
        .C1(n1949), .Y(n4199) );
  AOI211X1 U7553 ( .A0(n5917), .A1(n6475), .B0(n1966), .C0(n5793), .Y(n1965)
         );
  OAI222XL U7554 ( .A0(n1951), .A1(n5725), .B0(n1952), .B1(n5699), .C0(n6476), 
        .C1(n5750), .Y(n1966) );
  OAI222XL U7555 ( .A0(n1912), .A1(n6502), .B0(n1913), .B1(n5699), .C0(n6478), 
        .C1(n5750), .Y(n1927) );
  OAI222XL U7556 ( .A0(n1873), .A1(n5726), .B0(n1874), .B1(n5699), .C0(n6480), 
        .C1(n5750), .Y(n1888) );
  OAI222XL U7557 ( .A0(n1834), .A1(n5725), .B0(n1835), .B1(n5699), .C0(n6482), 
        .C1(n5750), .Y(n1849) );
  OAI222XL U7558 ( .A0(n6400), .A1(n5858), .B0(n1804), .B1(n1787), .C0(n269), 
        .C1(n1788), .Y(n4167) );
  AOI211X1 U7559 ( .A0(n5917), .A1(n6483), .B0(n1805), .C0(n5794), .Y(n1804)
         );
  OAI222XL U7560 ( .A0(n1790), .A1(n5726), .B0(n1791), .B1(n5699), .C0(n6484), 
        .C1(n5750), .Y(n1805) );
  OAI222XL U7561 ( .A0(n1745), .A1(n5725), .B0(n1746), .B1(n5699), .C0(n6486), 
        .C1(n5750), .Y(n1760) );
  OAI222XL U7562 ( .A0(n6402), .A1(n5858), .B0(n1715), .B1(n1698), .C0(n253), 
        .C1(n1699), .Y(n4151) );
  AOI211X1 U7563 ( .A0(N3375), .A1(n6487), .B0(n1716), .C0(n5794), .Y(n1715)
         );
  OAI222XL U7564 ( .A0(n1701), .A1(n6502), .B0(n1702), .B1(n5699), .C0(n6488), 
        .C1(n5750), .Y(n1716) );
  OAI222XL U7565 ( .A0(n6403), .A1(n5858), .B0(n1671), .B1(n1654), .C0(n245), 
        .C1(n1655), .Y(n4143) );
  AOI211X1 U7566 ( .A0(n5917), .A1(n6489), .B0(n1672), .C0(n5794), .Y(n1671)
         );
  OAI222XL U7567 ( .A0(n1657), .A1(n5726), .B0(n1658), .B1(n5699), .C0(n6490), 
        .C1(n5750), .Y(n1672) );
  OAI222XL U7568 ( .A0(n6404), .A1(n5858), .B0(n1627), .B1(n1610), .C0(n237), 
        .C1(n1611), .Y(n4135) );
  OAI222XL U7569 ( .A0(n1613), .A1(n5725), .B0(n1614), .B1(n5699), .C0(n6492), 
        .C1(n5750), .Y(n1628) );
  OAI222XL U7570 ( .A0(n6405), .A1(n5858), .B0(n1583), .B1(n1566), .C0(n229), 
        .C1(n1567), .Y(n4127) );
  AOI211X1 U7571 ( .A0(N3375), .A1(n6493), .B0(n1584), .C0(n5794), .Y(n1583)
         );
  OAI222XL U7572 ( .A0(n1569), .A1(n5724), .B0(n1570), .B1(n5699), .C0(n6494), 
        .C1(n5750), .Y(n1584) );
  OAI222XL U7573 ( .A0(n6406), .A1(n5857), .B0(n1539), .B1(n1522), .C0(n221), 
        .C1(n1523), .Y(n4119) );
  AOI211X1 U7574 ( .A0(n5917), .A1(n6495), .B0(n1540), .C0(n5794), .Y(n1539)
         );
  OAI222XL U7575 ( .A0(n1525), .A1(n5724), .B0(n1526), .B1(n5699), .C0(n6496), 
        .C1(n5750), .Y(n1540) );
  OAI222XL U7576 ( .A0(n6407), .A1(n5857), .B0(n1495), .B1(n1478), .C0(n213), 
        .C1(n1479), .Y(n4111) );
  OAI222XL U7577 ( .A0(n1481), .A1(n5724), .B0(n1482), .B1(n5701), .C0(n6498), 
        .C1(n5751), .Y(n1496) );
  OAI222XL U7578 ( .A0(n6347), .A1(n5863), .B0(n3945), .B1(n3929), .C0(n700), 
        .C1(n3930), .Y(n4598) );
  AOI211X1 U7579 ( .A0(n5921), .A1(n3931), .B0(n3946), .C0(n5860), .Y(n3945)
         );
  OAI222XL U7580 ( .A0(n3933), .A1(n5722), .B0(n3934), .B1(n5696), .C0(n6424), 
        .C1(n5747), .Y(n3946) );
  OAI222XL U7581 ( .A0(n6348), .A1(n5863), .B0(n3906), .B1(n3890), .C0(n692), 
        .C1(n3891), .Y(n4590) );
  AOI211X1 U7582 ( .A0(n5921), .A1(n3892), .B0(n3907), .C0(n5859), .Y(n3906)
         );
  OAI222XL U7583 ( .A0(n3894), .A1(n5722), .B0(n3895), .B1(n5697), .C0(n6425), 
        .C1(n5747), .Y(n3907) );
  OAI222XL U7584 ( .A0(n6349), .A1(n5863), .B0(n3867), .B1(n3851), .C0(n684), 
        .C1(n3852), .Y(n4582) );
  AOI211X1 U7585 ( .A0(n5921), .A1(n3853), .B0(n3868), .C0(n5861), .Y(n3867)
         );
  OAI222XL U7586 ( .A0(n3855), .A1(n5722), .B0(n3856), .B1(n5697), .C0(n6426), 
        .C1(n5748), .Y(n3868) );
  OAI222XL U7587 ( .A0(n6350), .A1(n5863), .B0(n3828), .B1(n3812), .C0(n676), 
        .C1(n3813), .Y(n4574) );
  AOI211X1 U7588 ( .A0(n5921), .A1(n3814), .B0(n3829), .C0(n5859), .Y(n3828)
         );
  OAI222XL U7589 ( .A0(n3816), .A1(n5722), .B0(n3817), .B1(n5697), .C0(n6427), 
        .C1(n5748), .Y(n3829) );
  OAI222XL U7590 ( .A0(n6351), .A1(n5863), .B0(n3789), .B1(n3773), .C0(n668), 
        .C1(n3774), .Y(n4566) );
  AOI211X1 U7591 ( .A0(n5921), .A1(n3775), .B0(n3790), .C0(n4698), .Y(n3789)
         );
  OAI222XL U7592 ( .A0(n3777), .A1(n5722), .B0(n3778), .B1(n5697), .C0(n6428), 
        .C1(n5748), .Y(n3790) );
  OAI222XL U7593 ( .A0(n6352), .A1(n5863), .B0(n3750), .B1(n3734), .C0(n660), 
        .C1(n3735), .Y(n4558) );
  AOI211X1 U7594 ( .A0(n5921), .A1(n3736), .B0(n3751), .C0(n5860), .Y(n3750)
         );
  OAI222XL U7595 ( .A0(n3738), .A1(n5722), .B0(n3739), .B1(n5697), .C0(n6429), 
        .C1(n5748), .Y(n3751) );
  OAI222XL U7596 ( .A0(n6353), .A1(n5863), .B0(n3706), .B1(n3690), .C0(n652), 
        .C1(n5670), .Y(n4550) );
  AOI211X1 U7597 ( .A0(n5921), .A1(n3692), .B0(n3707), .C0(n4698), .Y(n3706)
         );
  OAI222XL U7598 ( .A0(n3694), .A1(n5723), .B0(n3695), .B1(n5697), .C0(n6430), 
        .C1(n5748), .Y(n3707) );
  OAI222XL U7599 ( .A0(n6354), .A1(n5863), .B0(n3667), .B1(n3651), .C0(n644), 
        .C1(n3652), .Y(n4542) );
  AOI211X1 U7600 ( .A0(n5921), .A1(n3653), .B0(n3668), .C0(n5860), .Y(n3667)
         );
  OAI222XL U7601 ( .A0(n3655), .A1(n5722), .B0(n3656), .B1(n5697), .C0(n6431), 
        .C1(n5748), .Y(n3668) );
  OAI222XL U7602 ( .A0(n6355), .A1(n5863), .B0(n3628), .B1(n3612), .C0(n636), 
        .C1(n3613), .Y(n4534) );
  AOI211X1 U7603 ( .A0(n5921), .A1(n3614), .B0(n3629), .C0(n5859), .Y(n3628)
         );
  OAI222XL U7604 ( .A0(n3616), .A1(n5721), .B0(n3617), .B1(n5697), .C0(n6432), 
        .C1(n5748), .Y(n3629) );
  OAI222XL U7605 ( .A0(n6356), .A1(n5863), .B0(n3589), .B1(n3573), .C0(n628), 
        .C1(n3574), .Y(n4526) );
  AOI211X1 U7606 ( .A0(n5921), .A1(n3575), .B0(n3590), .C0(n4698), .Y(n3589)
         );
  OAI222XL U7607 ( .A0(n3577), .A1(n5722), .B0(n3578), .B1(n5697), .C0(n6433), 
        .C1(n5748), .Y(n3590) );
  OAI222XL U7608 ( .A0(n6357), .A1(n5863), .B0(n3550), .B1(n3534), .C0(n620), 
        .C1(n3535), .Y(n4518) );
  AOI211X1 U7609 ( .A0(n5921), .A1(n3536), .B0(n3551), .C0(n5860), .Y(n3550)
         );
  OAI222XL U7610 ( .A0(n3538), .A1(n5723), .B0(n3539), .B1(n5697), .C0(n6434), 
        .C1(n5748), .Y(n3551) );
  OAI222XL U7611 ( .A0(n6358), .A1(n5863), .B0(n3511), .B1(n3495), .C0(n612), 
        .C1(n3496), .Y(n4510) );
  AOI211X1 U7612 ( .A0(n5921), .A1(n3497), .B0(n3512), .C0(n4698), .Y(n3511)
         );
  OAI222XL U7613 ( .A0(n3499), .A1(n5721), .B0(n3500), .B1(n5697), .C0(n6435), 
        .C1(n5748), .Y(n3512) );
  OAI222XL U7614 ( .A0(n6359), .A1(n5865), .B0(n3472), .B1(n3456), .C0(n604), 
        .C1(n3457), .Y(n4502) );
  AOI211X1 U7615 ( .A0(n5921), .A1(n3458), .B0(n3473), .C0(n5859), .Y(n3472)
         );
  OAI222XL U7616 ( .A0(n3460), .A1(n5721), .B0(n3461), .B1(n5697), .C0(n6436), 
        .C1(n5748), .Y(n3473) );
  OAI222XL U7617 ( .A0(n6360), .A1(n5864), .B0(n3433), .B1(n3417), .C0(n596), 
        .C1(n3418), .Y(n4494) );
  AOI211X1 U7618 ( .A0(n5921), .A1(n3419), .B0(n3434), .C0(n5861), .Y(n3433)
         );
  OAI222XL U7619 ( .A0(n3421), .A1(n5721), .B0(n3422), .B1(n5697), .C0(n6437), 
        .C1(n5748), .Y(n3434) );
  OAI222XL U7620 ( .A0(n6361), .A1(n5863), .B0(n3389), .B1(n3373), .C0(n588), 
        .C1(n3374), .Y(n4486) );
  AOI211X1 U7621 ( .A0(n5921), .A1(n3375), .B0(n3390), .C0(n5859), .Y(n3389)
         );
  OAI222XL U7622 ( .A0(n3377), .A1(n5721), .B0(n3378), .B1(n5697), .C0(n6438), 
        .C1(n5748), .Y(n3390) );
  OAI222XL U7623 ( .A0(n6362), .A1(n5865), .B0(n3350), .B1(n3334), .C0(n580), 
        .C1(n3335), .Y(n4478) );
  AOI211X1 U7624 ( .A0(n5921), .A1(n3336), .B0(n3351), .C0(n5860), .Y(n3350)
         );
  OAI222XL U7625 ( .A0(n3338), .A1(n5721), .B0(n3339), .B1(n5697), .C0(n6439), 
        .C1(n5748), .Y(n3351) );
  OAI222XL U7626 ( .A0(n6363), .A1(n5864), .B0(n3311), .B1(n3295), .C0(n572), 
        .C1(n3296), .Y(n4470) );
  AOI211X1 U7627 ( .A0(n5921), .A1(n3297), .B0(n3312), .C0(n5860), .Y(n3311)
         );
  OAI222XL U7628 ( .A0(n3299), .A1(n5721), .B0(n3300), .B1(n5697), .C0(n6440), 
        .C1(n5748), .Y(n3312) );
  OAI222XL U7629 ( .A0(n6364), .A1(n5863), .B0(n3272), .B1(n3256), .C0(n564), 
        .C1(n3257), .Y(n4462) );
  AOI211X1 U7630 ( .A0(n5921), .A1(n3258), .B0(n3273), .C0(n4698), .Y(n3272)
         );
  OAI222XL U7631 ( .A0(n3260), .A1(n5721), .B0(n3261), .B1(n5697), .C0(n6441), 
        .C1(n5748), .Y(n3273) );
  OAI222XL U7632 ( .A0(n6365), .A1(n5865), .B0(n3233), .B1(n3217), .C0(n556), 
        .C1(n3218), .Y(n4454) );
  AOI211X1 U7633 ( .A0(n5921), .A1(n3219), .B0(n3234), .C0(n4698), .Y(n3233)
         );
  OAI222XL U7634 ( .A0(n3221), .A1(n5721), .B0(n3222), .B1(n5696), .C0(n6442), 
        .C1(n5748), .Y(n3234) );
  OAI222XL U7635 ( .A0(n6366), .A1(n5864), .B0(n3194), .B1(n3178), .C0(n548), 
        .C1(n3179), .Y(n4446) );
  AOI211X1 U7636 ( .A0(n5921), .A1(n3180), .B0(n3195), .C0(n5861), .Y(n3194)
         );
  OAI222XL U7637 ( .A0(n3182), .A1(n5721), .B0(n3183), .B1(n5695), .C0(n6443), 
        .C1(n5746), .Y(n3195) );
  OAI222XL U7638 ( .A0(n6367), .A1(n5864), .B0(n3155), .B1(n3139), .C0(n540), 
        .C1(n4674), .Y(n4438) );
  AOI211X1 U7639 ( .A0(n5921), .A1(n3141), .B0(n3156), .C0(n4698), .Y(n3155)
         );
  OAI222XL U7640 ( .A0(n3143), .A1(n5721), .B0(n3144), .B1(n5697), .C0(n6444), 
        .C1(n5748), .Y(n3156) );
  OAI222XL U7641 ( .A0(n6368), .A1(n5863), .B0(n3116), .B1(n3100), .C0(n532), 
        .C1(n3101), .Y(n4430) );
  AOI211X1 U7642 ( .A0(n5921), .A1(n3102), .B0(n3117), .C0(n5861), .Y(n3116)
         );
  OAI222XL U7643 ( .A0(n3104), .A1(n5721), .B0(n3105), .B1(n6036), .C0(n6445), 
        .C1(n5746), .Y(n3117) );
  OAI222XL U7644 ( .A0(n6369), .A1(n5865), .B0(n3072), .B1(n3056), .C0(n524), 
        .C1(n3057), .Y(n4422) );
  AOI211X1 U7645 ( .A0(n5921), .A1(n3058), .B0(n3073), .C0(n5861), .Y(n3072)
         );
  OAI222XL U7646 ( .A0(n3060), .A1(n5721), .B0(n3061), .B1(n5697), .C0(n6446), 
        .C1(n5748), .Y(n3073) );
  OAI222XL U7647 ( .A0(n6370), .A1(n5864), .B0(n3033), .B1(n3017), .C0(n516), 
        .C1(n3018), .Y(n4414) );
  AOI211X1 U7648 ( .A0(n5921), .A1(n3019), .B0(n3034), .C0(n5859), .Y(n3033)
         );
  OAI222XL U7649 ( .A0(n3021), .A1(n5722), .B0(n3022), .B1(n6422), .C0(n6447), 
        .C1(n5746), .Y(n3034) );
  OAI222XL U7650 ( .A0(n6371), .A1(n5864), .B0(n2994), .B1(n2978), .C0(n508), 
        .C1(n2979), .Y(n4406) );
  AOI211X1 U7651 ( .A0(n5921), .A1(n2980), .B0(n2995), .C0(n5860), .Y(n2994)
         );
  OAI222XL U7652 ( .A0(n2982), .A1(n5722), .B0(n2983), .B1(n5697), .C0(n6448), 
        .C1(n5748), .Y(n2995) );
  OAI222XL U7653 ( .A0(n6372), .A1(n5864), .B0(n2955), .B1(n2939), .C0(n500), 
        .C1(n4675), .Y(n4398) );
  AOI211X1 U7654 ( .A0(n5921), .A1(n2941), .B0(n2956), .C0(n5861), .Y(n2955)
         );
  OAI222XL U7655 ( .A0(n2943), .A1(n5722), .B0(n2944), .B1(n5696), .C0(n6449), 
        .C1(n5747), .Y(n2956) );
  OAI222XL U7656 ( .A0(n6373), .A1(n5864), .B0(n2916), .B1(n2900), .C0(n492), 
        .C1(n2901), .Y(n4390) );
  AOI211X1 U7657 ( .A0(n5921), .A1(n2902), .B0(n2917), .C0(n5859), .Y(n2916)
         );
  OAI222XL U7658 ( .A0(n2904), .A1(n5722), .B0(n2905), .B1(n6422), .C0(n6450), 
        .C1(n6508), .Y(n2917) );
  OAI222XL U7659 ( .A0(n6374), .A1(n5864), .B0(n2877), .B1(n2861), .C0(n484), 
        .C1(n2862), .Y(n4382) );
  AOI211X1 U7660 ( .A0(n5921), .A1(n2863), .B0(n2878), .C0(n5861), .Y(n2877)
         );
  OAI222XL U7661 ( .A0(n2865), .A1(n5722), .B0(n2866), .B1(n5697), .C0(n6451), 
        .C1(n5748), .Y(n2878) );
  OAI222XL U7662 ( .A0(n6375), .A1(n5864), .B0(n2838), .B1(n2822), .C0(n476), 
        .C1(n2823), .Y(n4374) );
  AOI211X1 U7663 ( .A0(n5921), .A1(n2824), .B0(n2839), .C0(n5860), .Y(n2838)
         );
  OAI222XL U7664 ( .A0(n2826), .A1(n5722), .B0(n2827), .B1(n6422), .C0(n6452), 
        .C1(n6508), .Y(n2839) );
  OAI222XL U7665 ( .A0(n6376), .A1(n5864), .B0(n2799), .B1(n2783), .C0(n468), 
        .C1(n2784), .Y(n4366) );
  AOI211X1 U7666 ( .A0(n5920), .A1(n2785), .B0(n2800), .C0(n4698), .Y(n2799)
         );
  OAI222XL U7667 ( .A0(n2787), .A1(n5722), .B0(n2788), .B1(n6422), .C0(n6453), 
        .C1(n6508), .Y(n2800) );
  OAI222XL U7668 ( .A0(n6377), .A1(n5864), .B0(n2755), .B1(n2739), .C0(n460), 
        .C1(n2740), .Y(n4358) );
  AOI211X1 U7669 ( .A0(n5920), .A1(n2741), .B0(n2756), .C0(n4698), .Y(n2755)
         );
  OAI222XL U7670 ( .A0(n2743), .A1(n5722), .B0(n2744), .B1(n6422), .C0(n6454), 
        .C1(n6508), .Y(n2756) );
  OAI222XL U7671 ( .A0(n6378), .A1(n5864), .B0(n2716), .B1(n2700), .C0(n452), 
        .C1(n2701), .Y(n4350) );
  AOI211X1 U7672 ( .A0(n5920), .A1(n2702), .B0(n2717), .C0(n4698), .Y(n2716)
         );
  OAI222XL U7673 ( .A0(n2704), .A1(n5722), .B0(n2705), .B1(n6422), .C0(n6455), 
        .C1(n6508), .Y(n2717) );
  OAI222XL U7674 ( .A0(n6379), .A1(n5864), .B0(n2677), .B1(n2661), .C0(n444), 
        .C1(n2662), .Y(n4342) );
  AOI211X1 U7675 ( .A0(n5920), .A1(n2663), .B0(n2678), .C0(n4698), .Y(n2677)
         );
  OAI222XL U7676 ( .A0(n2665), .A1(n5722), .B0(n2666), .B1(n5696), .C0(n6456), 
        .C1(n6508), .Y(n2678) );
  OAI222XL U7677 ( .A0(n6380), .A1(n5864), .B0(n2638), .B1(n2622), .C0(n436), 
        .C1(n2623), .Y(n4334) );
  AOI211X1 U7678 ( .A0(n5920), .A1(n2624), .B0(n2639), .C0(n4698), .Y(n2638)
         );
  OAI222XL U7679 ( .A0(n2626), .A1(n5722), .B0(n2627), .B1(n5696), .C0(n6457), 
        .C1(n5747), .Y(n2639) );
  OAI222XL U7680 ( .A0(n6381), .A1(n5864), .B0(n2599), .B1(n2583), .C0(n428), 
        .C1(n2584), .Y(n4326) );
  AOI211X1 U7681 ( .A0(n5920), .A1(n2585), .B0(n2600), .C0(n4698), .Y(n2599)
         );
  OAI222XL U7682 ( .A0(n2587), .A1(n5722), .B0(n2588), .B1(n5696), .C0(n6458), 
        .C1(n5747), .Y(n2600) );
  OAI222XL U7683 ( .A0(n6382), .A1(n5865), .B0(n2560), .B1(n2544), .C0(n420), 
        .C1(n2545), .Y(n4318) );
  AOI211X1 U7684 ( .A0(n5920), .A1(n2546), .B0(n2561), .C0(n5861), .Y(n2560)
         );
  OAI222XL U7685 ( .A0(n2548), .A1(n5721), .B0(n2549), .B1(n5696), .C0(n6459), 
        .C1(n5747), .Y(n2561) );
  OAI222XL U7686 ( .A0(n6383), .A1(n5865), .B0(n2521), .B1(n2505), .C0(n412), 
        .C1(n2506), .Y(n4310) );
  AOI211X1 U7687 ( .A0(n5920), .A1(n2507), .B0(n2522), .C0(n5859), .Y(n2521)
         );
  OAI222XL U7688 ( .A0(n2509), .A1(n5723), .B0(n2510), .B1(n5696), .C0(n6460), 
        .C1(n5747), .Y(n2522) );
  OAI222XL U7689 ( .A0(n6384), .A1(n5865), .B0(n2482), .B1(n2466), .C0(n404), 
        .C1(n2467), .Y(n4302) );
  AOI211X1 U7690 ( .A0(n5920), .A1(n2468), .B0(n2483), .C0(n4698), .Y(n2482)
         );
  OAI222XL U7691 ( .A0(n2470), .A1(n5721), .B0(n2471), .B1(n5696), .C0(n6461), 
        .C1(n5747), .Y(n2483) );
  OAI222XL U7692 ( .A0(n6385), .A1(n5865), .B0(n2438), .B1(n2422), .C0(n396), 
        .C1(n2423), .Y(n4294) );
  AOI211X1 U7693 ( .A0(n5920), .A1(n2424), .B0(n2439), .C0(n4698), .Y(n2438)
         );
  OAI222XL U7694 ( .A0(n2426), .A1(n5723), .B0(n2427), .B1(n5696), .C0(n6462), 
        .C1(n5747), .Y(n2439) );
  OAI222XL U7695 ( .A0(n6386), .A1(n5865), .B0(n2399), .B1(n2383), .C0(n388), 
        .C1(n2384), .Y(n4286) );
  AOI211X1 U7696 ( .A0(n5920), .A1(n2385), .B0(n2400), .C0(n5860), .Y(n2399)
         );
  OAI222XL U7697 ( .A0(n2387), .A1(n5721), .B0(n2388), .B1(n5696), .C0(n6463), 
        .C1(n5747), .Y(n2400) );
  OAI222XL U7698 ( .A0(n6387), .A1(n5865), .B0(n2360), .B1(n2344), .C0(n380), 
        .C1(n2345), .Y(n4278) );
  AOI211X1 U7699 ( .A0(n5920), .A1(n2346), .B0(n2361), .C0(n5861), .Y(n2360)
         );
  OAI222XL U7700 ( .A0(n2348), .A1(n5723), .B0(n2349), .B1(n5696), .C0(n6464), 
        .C1(n5747), .Y(n2361) );
  OAI222XL U7701 ( .A0(n6388), .A1(n5865), .B0(n2321), .B1(n2305), .C0(n372), 
        .C1(n2306), .Y(n4270) );
  AOI211X1 U7702 ( .A0(n5920), .A1(n2307), .B0(n2322), .C0(n5859), .Y(n2321)
         );
  OAI222XL U7703 ( .A0(n2309), .A1(n5721), .B0(n2310), .B1(n5696), .C0(n6465), 
        .C1(n5747), .Y(n2322) );
  OAI222XL U7704 ( .A0(n6389), .A1(n5865), .B0(n2282), .B1(n2266), .C0(n364), 
        .C1(n2267), .Y(n4262) );
  AOI211X1 U7705 ( .A0(n5920), .A1(n2268), .B0(n2283), .C0(n4698), .Y(n2282)
         );
  OAI222XL U7706 ( .A0(n2270), .A1(n5721), .B0(n2271), .B1(n5696), .C0(n6466), 
        .C1(n5747), .Y(n2283) );
  OAI222XL U7707 ( .A0(n6390), .A1(n5865), .B0(n2243), .B1(n2227), .C0(n356), 
        .C1(n2228), .Y(n4254) );
  AOI211X1 U7708 ( .A0(n5920), .A1(n2229), .B0(n2244), .C0(n4698), .Y(n2243)
         );
  OAI222XL U7709 ( .A0(n2231), .A1(n5723), .B0(n2232), .B1(n5696), .C0(n6467), 
        .C1(n5747), .Y(n2244) );
  OAI222XL U7710 ( .A0(n6391), .A1(n5865), .B0(n2204), .B1(n2188), .C0(n348), 
        .C1(n2189), .Y(n4246) );
  AOI211X1 U7711 ( .A0(n5920), .A1(n2190), .B0(n2205), .C0(n5860), .Y(n2204)
         );
  OAI222XL U7712 ( .A0(n2192), .A1(n5723), .B0(n2193), .B1(n5696), .C0(n6468), 
        .C1(n5747), .Y(n2205) );
  OAI222XL U7713 ( .A0(n6392), .A1(n5865), .B0(n2165), .B1(n2149), .C0(n340), 
        .C1(n2150), .Y(n4238) );
  AOI211X1 U7714 ( .A0(n5920), .A1(n2151), .B0(n2166), .C0(n5861), .Y(n2165)
         );
  OAI222XL U7715 ( .A0(n2153), .A1(n5721), .B0(n2154), .B1(n5696), .C0(n6469), 
        .C1(n5747), .Y(n2166) );
  OAI222XL U7716 ( .A0(n6393), .A1(n5865), .B0(n2121), .B1(n2105), .C0(n332), 
        .C1(n2106), .Y(n4230) );
  AOI211X1 U7717 ( .A0(n5920), .A1(n2107), .B0(n2122), .C0(n5859), .Y(n2121)
         );
  OAI222XL U7718 ( .A0(n2109), .A1(n5723), .B0(n2110), .B1(n5696), .C0(n6470), 
        .C1(n5747), .Y(n2122) );
  OAI222XL U7719 ( .A0(n6394), .A1(n5864), .B0(n2082), .B1(n2066), .C0(n324), 
        .C1(n2067), .Y(n4222) );
  AOI211X1 U7720 ( .A0(n5920), .A1(n2068), .B0(n2083), .C0(n4698), .Y(n2082)
         );
  OAI222XL U7721 ( .A0(n2070), .A1(n5723), .B0(n2071), .B1(n5696), .C0(n6471), 
        .C1(n5747), .Y(n2083) );
  OAI222XL U7722 ( .A0(n6395), .A1(n5863), .B0(n2043), .B1(n2027), .C0(n316), 
        .C1(n2028), .Y(n4214) );
  AOI211X1 U7723 ( .A0(n5920), .A1(n2029), .B0(n2044), .C0(n4698), .Y(n2043)
         );
  OAI222XL U7724 ( .A0(n2031), .A1(n5723), .B0(n2032), .B1(n5695), .C0(n6472), 
        .C1(n5747), .Y(n2044) );
  OAI222XL U7725 ( .A0(n1990), .A1(n5723), .B0(n1991), .B1(n5695), .C0(n6474), 
        .C1(n5746), .Y(n2003) );
  OAI222XL U7726 ( .A0(n6397), .A1(n5865), .B0(n1963), .B1(n1948), .C0(n300), 
        .C1(n1949), .Y(n4198) );
  AOI211X1 U7727 ( .A0(n5920), .A1(n6475), .B0(n1964), .C0(n5860), .Y(n1963)
         );
  OAI222XL U7728 ( .A0(n1951), .A1(n5723), .B0(n1952), .B1(n5695), .C0(n6476), 
        .C1(n5746), .Y(n1964) );
  OAI222XL U7729 ( .A0(n6398), .A1(n5863), .B0(n1924), .B1(n1909), .C0(n292), 
        .C1(n1910), .Y(n4190) );
  AOI211X1 U7730 ( .A0(n5920), .A1(n6477), .B0(n1925), .C0(n5861), .Y(n1924)
         );
  OAI222XL U7731 ( .A0(n1912), .A1(n5723), .B0(n1913), .B1(n5695), .C0(n6478), 
        .C1(n5746), .Y(n1925) );
  OAI222XL U7732 ( .A0(n4832), .A1(n5865), .B0(n1885), .B1(n1870), .C0(n284), 
        .C1(n1871), .Y(n4182) );
  AOI211X1 U7733 ( .A0(n5920), .A1(n6479), .B0(n1886), .C0(n5859), .Y(n1885)
         );
  OAI222XL U7734 ( .A0(n1873), .A1(n5723), .B0(n1874), .B1(n5695), .C0(n6480), 
        .C1(n5746), .Y(n1886) );
  OAI222XL U7735 ( .A0(n1834), .A1(n5723), .B0(n1835), .B1(n5695), .C0(n6482), 
        .C1(n5746), .Y(n1847) );
  OAI222XL U7736 ( .A0(n6400), .A1(n5863), .B0(n1802), .B1(n1787), .C0(n268), 
        .C1(n1788), .Y(n4166) );
  AOI211X1 U7737 ( .A0(n5920), .A1(n6483), .B0(n1803), .C0(n4698), .Y(n1802)
         );
  OAI222XL U7738 ( .A0(n1790), .A1(n5723), .B0(n1791), .B1(n5695), .C0(n6484), 
        .C1(n5746), .Y(n1803) );
  OAI222XL U7739 ( .A0(n6401), .A1(n5864), .B0(n1757), .B1(n1742), .C0(n260), 
        .C1(n1743), .Y(n4158) );
  AOI211X1 U7740 ( .A0(n5920), .A1(n6485), .B0(n1758), .C0(n5860), .Y(n1757)
         );
  OAI222XL U7741 ( .A0(n1745), .A1(n5723), .B0(n1746), .B1(n5695), .C0(n6486), 
        .C1(n5746), .Y(n1758) );
  OAI222XL U7742 ( .A0(n6402), .A1(n5863), .B0(n1713), .B1(n1698), .C0(n252), 
        .C1(n1699), .Y(n4150) );
  AOI211X1 U7743 ( .A0(n5920), .A1(n6487), .B0(n1714), .C0(n5859), .Y(n1713)
         );
  OAI222XL U7744 ( .A0(n1701), .A1(n5723), .B0(n1702), .B1(n5695), .C0(n6488), 
        .C1(n5746), .Y(n1714) );
  OAI222XL U7745 ( .A0(n6403), .A1(n5865), .B0(n1669), .B1(n1654), .C0(n244), 
        .C1(n1655), .Y(n4142) );
  AOI211X1 U7746 ( .A0(n5920), .A1(n6489), .B0(n1670), .C0(n4698), .Y(n1669)
         );
  OAI222XL U7747 ( .A0(n1657), .A1(n5723), .B0(n1658), .B1(n5695), .C0(n6490), 
        .C1(n5746), .Y(n1670) );
  OAI222XL U7748 ( .A0(n6404), .A1(n5865), .B0(n1625), .B1(n1610), .C0(n236), 
        .C1(n1611), .Y(n4134) );
  AOI211X1 U7749 ( .A0(n5920), .A1(n6491), .B0(n1626), .C0(n5860), .Y(n1625)
         );
  OAI222XL U7750 ( .A0(n1613), .A1(n5723), .B0(n1614), .B1(n5695), .C0(n6492), 
        .C1(n5746), .Y(n1626) );
  OAI222XL U7751 ( .A0(n6405), .A1(n5864), .B0(n1581), .B1(n1566), .C0(n228), 
        .C1(n1567), .Y(n4126) );
  AOI211X1 U7752 ( .A0(n5920), .A1(n6493), .B0(n1582), .C0(n4698), .Y(n1581)
         );
  OAI222XL U7753 ( .A0(n1569), .A1(n5721), .B0(n1570), .B1(n5695), .C0(n6494), 
        .C1(n5746), .Y(n1582) );
  OAI222XL U7754 ( .A0(n6406), .A1(n5863), .B0(n1537), .B1(n1522), .C0(n220), 
        .C1(n1523), .Y(n4118) );
  AOI211X1 U7755 ( .A0(n5920), .A1(n6495), .B0(n1538), .C0(n5861), .Y(n1537)
         );
  OAI222XL U7756 ( .A0(n1525), .A1(n5721), .B0(n1526), .B1(n5695), .C0(n6496), 
        .C1(n5746), .Y(n1538) );
  OAI222XL U7757 ( .A0(n6407), .A1(n5865), .B0(n1493), .B1(n1478), .C0(n212), 
        .C1(n1479), .Y(n4110) );
  AOI211X1 U7758 ( .A0(n5921), .A1(n6497), .B0(n1494), .C0(n4698), .Y(n1493)
         );
  OAI222XL U7759 ( .A0(n1481), .A1(n5723), .B0(n1482), .B1(n5696), .C0(n6498), 
        .C1(n5747), .Y(n1494) );
  OAI222XL U7760 ( .A0(n6347), .A1(n5872), .B0(n3943), .B1(n3929), .C0(n699), 
        .C1(n3930), .Y(n4597) );
  OAI222XL U7761 ( .A0(n3933), .A1(n5718), .B0(n3934), .B1(n5692), .C0(n6424), 
        .C1(n5744), .Y(n3944) );
  OAI222XL U7762 ( .A0(n6348), .A1(n5872), .B0(n3904), .B1(n3890), .C0(n691), 
        .C1(n3891), .Y(n4589) );
  OAI222XL U7763 ( .A0(n3894), .A1(n5718), .B0(n3895), .B1(n5694), .C0(n6425), 
        .C1(n5744), .Y(n3905) );
  OAI222XL U7764 ( .A0(n6349), .A1(n5872), .B0(n3865), .B1(n3851), .C0(n683), 
        .C1(n3852), .Y(n4581) );
  OAI222XL U7765 ( .A0(n3855), .A1(n5718), .B0(n3856), .B1(n5694), .C0(n6426), 
        .C1(n5743), .Y(n3866) );
  OAI222XL U7766 ( .A0(n6350), .A1(n5872), .B0(n3826), .B1(n3812), .C0(n675), 
        .C1(n3813), .Y(n4573) );
  OAI222XL U7767 ( .A0(n3816), .A1(n5718), .B0(n3817), .B1(n5694), .C0(n6427), 
        .C1(n5743), .Y(n3827) );
  OAI222XL U7768 ( .A0(n6351), .A1(n5872), .B0(n3787), .B1(n3773), .C0(n667), 
        .C1(n3774), .Y(n4565) );
  OAI222XL U7769 ( .A0(n3777), .A1(n5718), .B0(n3778), .B1(n5694), .C0(n6428), 
        .C1(n5743), .Y(n3788) );
  OAI222XL U7770 ( .A0(n6352), .A1(n5872), .B0(n3748), .B1(n3734), .C0(n659), 
        .C1(n3735), .Y(n4557) );
  OAI222XL U7771 ( .A0(n3738), .A1(n5718), .B0(n3739), .B1(n5694), .C0(n6429), 
        .C1(n6507), .Y(n3749) );
  OAI222XL U7772 ( .A0(n6353), .A1(n5872), .B0(n3704), .B1(n3690), .C0(n651), 
        .C1(n5670), .Y(n4549) );
  OAI222XL U7773 ( .A0(n3694), .A1(n5718), .B0(n3695), .B1(n5694), .C0(n6430), 
        .C1(n6507), .Y(n3705) );
  OAI222XL U7774 ( .A0(n6354), .A1(n5872), .B0(n3665), .B1(n3651), .C0(n643), 
        .C1(n3652), .Y(n4541) );
  OAI222XL U7775 ( .A0(n3655), .A1(n5718), .B0(n3656), .B1(n5694), .C0(n6431), 
        .C1(n6507), .Y(n3666) );
  OAI222XL U7776 ( .A0(n6355), .A1(n5872), .B0(n3626), .B1(n3612), .C0(n635), 
        .C1(n3613), .Y(n4533) );
  OAI222XL U7777 ( .A0(n3616), .A1(n5718), .B0(n3617), .B1(n5694), .C0(n6432), 
        .C1(n6507), .Y(n3627) );
  OAI222XL U7778 ( .A0(n6356), .A1(n5872), .B0(n3587), .B1(n3573), .C0(n627), 
        .C1(n3574), .Y(n4525) );
  OAI222XL U7779 ( .A0(n3577), .A1(n5718), .B0(n3578), .B1(n5694), .C0(n6433), 
        .C1(n6507), .Y(n3588) );
  OAI222XL U7780 ( .A0(n6357), .A1(n5872), .B0(n3548), .B1(n3534), .C0(n619), 
        .C1(n3535), .Y(n4517) );
  OAI222XL U7781 ( .A0(n3538), .A1(n5718), .B0(n3539), .B1(n5694), .C0(n6434), 
        .C1(n5743), .Y(n3549) );
  OAI222XL U7782 ( .A0(n6358), .A1(n5872), .B0(n3509), .B1(n3495), .C0(n611), 
        .C1(n3496), .Y(n4509) );
  OAI222XL U7783 ( .A0(n3499), .A1(n5719), .B0(n3500), .B1(n5694), .C0(n6435), 
        .C1(n5745), .Y(n3510) );
  OAI222XL U7784 ( .A0(n6359), .A1(n5874), .B0(n3470), .B1(n3456), .C0(n603), 
        .C1(n3457), .Y(n4501) );
  OAI222XL U7785 ( .A0(n3460), .A1(n5719), .B0(n3461), .B1(n5694), .C0(n6436), 
        .C1(n5744), .Y(n3471) );
  OAI222XL U7786 ( .A0(n6360), .A1(n5873), .B0(n3431), .B1(n3417), .C0(n595), 
        .C1(n3418), .Y(n4493) );
  OAI222XL U7787 ( .A0(n3421), .A1(n5719), .B0(n3422), .B1(n5694), .C0(n6437), 
        .C1(n5744), .Y(n3432) );
  OAI222XL U7788 ( .A0(n6361), .A1(n5875), .B0(n3387), .B1(n3373), .C0(n587), 
        .C1(n3374), .Y(n4485) );
  OAI222XL U7789 ( .A0(n3377), .A1(n5719), .B0(n3378), .B1(n5694), .C0(n6438), 
        .C1(n5745), .Y(n3388) );
  OAI222XL U7790 ( .A0(n6362), .A1(n5875), .B0(n3348), .B1(n3334), .C0(n579), 
        .C1(n3335), .Y(n4477) );
  OAI222XL U7791 ( .A0(n3338), .A1(n5719), .B0(n3339), .B1(n5694), .C0(n6439), 
        .C1(n5745), .Y(n3349) );
  OAI222XL U7792 ( .A0(n6363), .A1(n5872), .B0(n3309), .B1(n3295), .C0(n571), 
        .C1(n3296), .Y(n4469) );
  OAI222XL U7793 ( .A0(n3299), .A1(n5719), .B0(n3300), .B1(n5694), .C0(n6440), 
        .C1(n5745), .Y(n3310) );
  OAI222XL U7794 ( .A0(n6364), .A1(n5872), .B0(n3270), .B1(n3256), .C0(n563), 
        .C1(n3257), .Y(n4461) );
  OAI222XL U7795 ( .A0(n3260), .A1(n5719), .B0(n3261), .B1(n5693), .C0(n6441), 
        .C1(n5745), .Y(n3271) );
  OAI222XL U7796 ( .A0(n6365), .A1(n5874), .B0(n3231), .B1(n3217), .C0(n555), 
        .C1(n3218), .Y(n4453) );
  OAI222XL U7797 ( .A0(n3221), .A1(n5719), .B0(n3222), .B1(n5693), .C0(n6442), 
        .C1(n5745), .Y(n3232) );
  OAI222XL U7798 ( .A0(n6366), .A1(n5874), .B0(n3192), .B1(n3178), .C0(n547), 
        .C1(n3179), .Y(n4445) );
  OAI222XL U7799 ( .A0(n3182), .A1(n5719), .B0(n3183), .B1(n5693), .C0(n6443), 
        .C1(n5745), .Y(n3193) );
  OAI222XL U7800 ( .A0(n6367), .A1(n5873), .B0(n3153), .B1(n3139), .C0(n539), 
        .C1(n4674), .Y(n4437) );
  OAI222XL U7801 ( .A0(n3143), .A1(n5719), .B0(n3144), .B1(n5693), .C0(n6444), 
        .C1(n5745), .Y(n3154) );
  OAI222XL U7802 ( .A0(n6368), .A1(n5873), .B0(n3114), .B1(n3100), .C0(n531), 
        .C1(n3101), .Y(n4429) );
  OAI222XL U7803 ( .A0(n3104), .A1(n5719), .B0(n3105), .B1(n5693), .C0(n6445), 
        .C1(n5745), .Y(n3115) );
  OAI222XL U7804 ( .A0(n6369), .A1(n5873), .B0(n3070), .B1(n3056), .C0(n523), 
        .C1(n3057), .Y(n4421) );
  OAI222XL U7805 ( .A0(n3060), .A1(n5719), .B0(n3061), .B1(n5693), .C0(n6446), 
        .C1(n5745), .Y(n3071) );
  OAI222XL U7806 ( .A0(n6370), .A1(n5873), .B0(n3031), .B1(n3017), .C0(n515), 
        .C1(n3018), .Y(n4413) );
  OAI222XL U7807 ( .A0(n3021), .A1(n5720), .B0(n3022), .B1(n5693), .C0(n6447), 
        .C1(n5745), .Y(n3032) );
  OAI222XL U7808 ( .A0(n6371), .A1(n5873), .B0(n2992), .B1(n2978), .C0(n507), 
        .C1(n2979), .Y(n4405) );
  OAI222XL U7809 ( .A0(n2982), .A1(n5720), .B0(n2983), .B1(n5693), .C0(n6448), 
        .C1(n5745), .Y(n2993) );
  OAI222XL U7810 ( .A0(n6372), .A1(n5873), .B0(n2953), .B1(n2939), .C0(n499), 
        .C1(n4675), .Y(n4397) );
  OAI222XL U7811 ( .A0(n2943), .A1(n5720), .B0(n2944), .B1(n5693), .C0(n6449), 
        .C1(n5745), .Y(n2954) );
  OAI222XL U7812 ( .A0(n6373), .A1(n5873), .B0(n2914), .B1(n2900), .C0(n491), 
        .C1(n2901), .Y(n4389) );
  OAI222XL U7813 ( .A0(n2904), .A1(n5720), .B0(n2905), .B1(n5693), .C0(n6450), 
        .C1(n5745), .Y(n2915) );
  OAI222XL U7814 ( .A0(n6374), .A1(n5873), .B0(n2875), .B1(n2861), .C0(n483), 
        .C1(n2862), .Y(n4381) );
  OAI222XL U7815 ( .A0(n2865), .A1(n5720), .B0(n2866), .B1(n5693), .C0(n6451), 
        .C1(n5745), .Y(n2876) );
  OAI222XL U7816 ( .A0(n6375), .A1(n5873), .B0(n2836), .B1(n2822), .C0(n475), 
        .C1(n2823), .Y(n4373) );
  OAI222XL U7817 ( .A0(n2826), .A1(n5720), .B0(n2827), .B1(n5693), .C0(n6452), 
        .C1(n5745), .Y(n2837) );
  OAI222XL U7818 ( .A0(n6376), .A1(n5873), .B0(n2797), .B1(n2783), .C0(n467), 
        .C1(n2784), .Y(n4365) );
  AOI211X1 U7819 ( .A0(n5925), .A1(n2785), .B0(n2798), .C0(n5867), .Y(n2797)
         );
  OAI222XL U7820 ( .A0(n2787), .A1(n5720), .B0(n2788), .B1(n5693), .C0(n6453), 
        .C1(n5745), .Y(n2798) );
  OAI222XL U7821 ( .A0(n6377), .A1(n5873), .B0(n2753), .B1(n2739), .C0(n459), 
        .C1(n2740), .Y(n4357) );
  AOI211X1 U7822 ( .A0(n5925), .A1(n2741), .B0(n2754), .C0(n5867), .Y(n2753)
         );
  OAI222XL U7823 ( .A0(n2743), .A1(n5720), .B0(n2744), .B1(n5693), .C0(n6454), 
        .C1(n5745), .Y(n2754) );
  OAI222XL U7824 ( .A0(n6378), .A1(n5873), .B0(n2714), .B1(n2700), .C0(n451), 
        .C1(n2701), .Y(n4349) );
  AOI211X1 U7825 ( .A0(n5925), .A1(n2702), .B0(n2715), .C0(n5867), .Y(n2714)
         );
  OAI222XL U7826 ( .A0(n2704), .A1(n5720), .B0(n2705), .B1(n5693), .C0(n6455), 
        .C1(n5745), .Y(n2715) );
  OAI222XL U7827 ( .A0(n6379), .A1(n5873), .B0(n2675), .B1(n2661), .C0(n443), 
        .C1(n2662), .Y(n4341) );
  AOI211X1 U7828 ( .A0(n5925), .A1(n2663), .B0(n2676), .C0(n5867), .Y(n2675)
         );
  OAI222XL U7829 ( .A0(n2665), .A1(n5720), .B0(n2666), .B1(n5692), .C0(n6456), 
        .C1(n5745), .Y(n2676) );
  OAI222XL U7830 ( .A0(n6380), .A1(n5873), .B0(n2636), .B1(n2622), .C0(n435), 
        .C1(n2623), .Y(n4333) );
  AOI211X1 U7831 ( .A0(n5925), .A1(n2624), .B0(n2637), .C0(n5867), .Y(n2636)
         );
  OAI222XL U7832 ( .A0(n2626), .A1(n5720), .B0(n2627), .B1(n5692), .C0(n6457), 
        .C1(n5744), .Y(n2637) );
  OAI222XL U7833 ( .A0(n6381), .A1(n5873), .B0(n2597), .B1(n2583), .C0(n427), 
        .C1(n2584), .Y(n4325) );
  AOI211X1 U7834 ( .A0(n5925), .A1(n2585), .B0(n2598), .C0(n5867), .Y(n2597)
         );
  OAI222XL U7835 ( .A0(n2587), .A1(n5720), .B0(n2588), .B1(n5692), .C0(n6458), 
        .C1(n5744), .Y(n2598) );
  OAI222XL U7836 ( .A0(n6382), .A1(n5874), .B0(n2558), .B1(n2544), .C0(n419), 
        .C1(n2545), .Y(n4317) );
  AOI211X1 U7837 ( .A0(n5925), .A1(n2546), .B0(n2559), .C0(n5867), .Y(n2558)
         );
  OAI222XL U7838 ( .A0(n2548), .A1(n5720), .B0(n2549), .B1(n5692), .C0(n6459), 
        .C1(n5744), .Y(n2559) );
  OAI222XL U7839 ( .A0(n6383), .A1(n5874), .B0(n2519), .B1(n2505), .C0(n411), 
        .C1(n2506), .Y(n4309) );
  AOI211X1 U7840 ( .A0(n5925), .A1(n2507), .B0(n2520), .C0(n5867), .Y(n2519)
         );
  OAI222XL U7841 ( .A0(n2509), .A1(n5719), .B0(n2510), .B1(n5692), .C0(n6460), 
        .C1(n5744), .Y(n2520) );
  OAI222XL U7842 ( .A0(n6384), .A1(n5874), .B0(n2480), .B1(n2466), .C0(n403), 
        .C1(n2467), .Y(n4301) );
  AOI211X1 U7843 ( .A0(n5925), .A1(n2468), .B0(n2481), .C0(n5867), .Y(n2480)
         );
  OAI222XL U7844 ( .A0(n2470), .A1(n5720), .B0(n2471), .B1(n5692), .C0(n6461), 
        .C1(n5744), .Y(n2481) );
  OAI222XL U7845 ( .A0(n6385), .A1(n5874), .B0(n2436), .B1(n2422), .C0(n395), 
        .C1(n2423), .Y(n4293) );
  AOI211X1 U7846 ( .A0(n5925), .A1(n2424), .B0(n2437), .C0(n5868), .Y(n2436)
         );
  OAI222XL U7847 ( .A0(n2426), .A1(n5719), .B0(n2427), .B1(n5692), .C0(n6462), 
        .C1(n5744), .Y(n2437) );
  OAI222XL U7848 ( .A0(n6386), .A1(n5874), .B0(n2397), .B1(n2383), .C0(n387), 
        .C1(n2384), .Y(n4285) );
  AOI211X1 U7849 ( .A0(n5925), .A1(n2385), .B0(n2398), .C0(n5868), .Y(n2397)
         );
  OAI222XL U7850 ( .A0(n2387), .A1(n5720), .B0(n2388), .B1(n5692), .C0(n6463), 
        .C1(n5744), .Y(n2398) );
  OAI222XL U7851 ( .A0(n6387), .A1(n5874), .B0(n2358), .B1(n2344), .C0(n379), 
        .C1(n2345), .Y(n4277) );
  AOI211X1 U7852 ( .A0(n5925), .A1(n2346), .B0(n2359), .C0(n5868), .Y(n2358)
         );
  OAI222XL U7853 ( .A0(n2348), .A1(n5719), .B0(n2349), .B1(n5692), .C0(n6464), 
        .C1(n5744), .Y(n2359) );
  OAI222XL U7854 ( .A0(n6388), .A1(n5874), .B0(n2319), .B1(n2305), .C0(n371), 
        .C1(n2306), .Y(n4269) );
  AOI211X1 U7855 ( .A0(n5925), .A1(n2307), .B0(n2320), .C0(n5868), .Y(n2319)
         );
  OAI222XL U7856 ( .A0(n2309), .A1(n5720), .B0(n2310), .B1(n5692), .C0(n6465), 
        .C1(n5744), .Y(n2320) );
  OAI222XL U7857 ( .A0(n6389), .A1(n5874), .B0(n2280), .B1(n2266), .C0(n363), 
        .C1(n2267), .Y(n4261) );
  AOI211X1 U7858 ( .A0(n5925), .A1(n2268), .B0(n2281), .C0(n5868), .Y(n2280)
         );
  OAI222XL U7859 ( .A0(n2270), .A1(n5719), .B0(n2271), .B1(n5692), .C0(n6466), 
        .C1(n5744), .Y(n2281) );
  OAI222XL U7860 ( .A0(n6390), .A1(n5874), .B0(n2241), .B1(n2227), .C0(n355), 
        .C1(n2228), .Y(n4253) );
  AOI211X1 U7861 ( .A0(n5925), .A1(n2229), .B0(n2242), .C0(n5868), .Y(n2241)
         );
  OAI222XL U7862 ( .A0(n2231), .A1(n5720), .B0(n2232), .B1(n5692), .C0(n6467), 
        .C1(n5744), .Y(n2242) );
  OAI222XL U7863 ( .A0(n6391), .A1(n5874), .B0(n2202), .B1(n2188), .C0(n347), 
        .C1(n2189), .Y(n4245) );
  AOI211X1 U7864 ( .A0(n5925), .A1(n2190), .B0(n2203), .C0(n5868), .Y(n2202)
         );
  OAI222XL U7865 ( .A0(n2192), .A1(n5718), .B0(n2193), .B1(n5692), .C0(n6468), 
        .C1(n5744), .Y(n2203) );
  OAI222XL U7866 ( .A0(n6392), .A1(n5874), .B0(n2163), .B1(n2149), .C0(n339), 
        .C1(n2150), .Y(n4237) );
  AOI211X1 U7867 ( .A0(n5925), .A1(n2151), .B0(n2164), .C0(n5868), .Y(n2163)
         );
  OAI222XL U7868 ( .A0(n2153), .A1(n6501), .B0(n2154), .B1(n5692), .C0(n6469), 
        .C1(n5744), .Y(n2164) );
  OAI222XL U7869 ( .A0(n6393), .A1(n5874), .B0(n2119), .B1(n2105), .C0(n331), 
        .C1(n2106), .Y(n4229) );
  AOI211X1 U7870 ( .A0(n5925), .A1(n2107), .B0(n2120), .C0(n5868), .Y(n2119)
         );
  OAI222XL U7871 ( .A0(n2109), .A1(n4808), .B0(n2110), .B1(n5692), .C0(n6470), 
        .C1(n5744), .Y(n2120) );
  OAI222XL U7872 ( .A0(n6394), .A1(n5875), .B0(n2080), .B1(n2066), .C0(n323), 
        .C1(n2067), .Y(n4221) );
  AOI211X1 U7873 ( .A0(n5925), .A1(n2068), .B0(n2081), .C0(n5868), .Y(n2080)
         );
  OAI222XL U7874 ( .A0(n2070), .A1(n5719), .B0(n2071), .B1(n5692), .C0(n6471), 
        .C1(n5744), .Y(n2081) );
  OAI222XL U7875 ( .A0(n6395), .A1(n5875), .B0(n2041), .B1(n2027), .C0(n315), 
        .C1(n2028), .Y(n4213) );
  AOI211X1 U7876 ( .A0(n5925), .A1(n2029), .B0(n2042), .C0(n5868), .Y(n2041)
         );
  OAI222XL U7877 ( .A0(n2031), .A1(n5719), .B0(n2032), .B1(n5691), .C0(n6472), 
        .C1(n5744), .Y(n2042) );
  OAI222XL U7878 ( .A0(n6396), .A1(n5875), .B0(n2000), .B1(n1987), .C0(n307), 
        .C1(n1988), .Y(n4205) );
  AOI211X1 U7879 ( .A0(n5925), .A1(n6473), .B0(n2001), .C0(n5868), .Y(n2000)
         );
  OAI222XL U7880 ( .A0(n1990), .A1(n6501), .B0(n1991), .B1(n5691), .C0(n6474), 
        .C1(n5743), .Y(n2001) );
  OAI222XL U7881 ( .A0(n6397), .A1(n5875), .B0(n1961), .B1(n1948), .C0(n299), 
        .C1(n1949), .Y(n4197) );
  AOI211X1 U7882 ( .A0(n5925), .A1(n6475), .B0(n1962), .C0(n5868), .Y(n1961)
         );
  OAI222XL U7883 ( .A0(n1951), .A1(n5720), .B0(n1952), .B1(n5691), .C0(n6476), 
        .C1(n5743), .Y(n1962) );
  OAI222XL U7884 ( .A0(n6398), .A1(n5875), .B0(n1922), .B1(n1909), .C0(n291), 
        .C1(n1910), .Y(n4189) );
  AOI211X1 U7885 ( .A0(n5925), .A1(n6477), .B0(n1923), .C0(n5869), .Y(n1922)
         );
  OAI222XL U7886 ( .A0(n1912), .A1(n5720), .B0(n1913), .B1(n5691), .C0(n6478), 
        .C1(n5743), .Y(n1923) );
  OAI222XL U7887 ( .A0(n4832), .A1(n5875), .B0(n1883), .B1(n1870), .C0(n283), 
        .C1(n1871), .Y(n4181) );
  AOI211X1 U7888 ( .A0(n5925), .A1(n6479), .B0(n1884), .C0(n5869), .Y(n1883)
         );
  OAI222XL U7889 ( .A0(n1873), .A1(n6501), .B0(n1874), .B1(n5691), .C0(n6480), 
        .C1(n5743), .Y(n1884) );
  AOI211X1 U7890 ( .A0(n5925), .A1(n6481), .B0(n1845), .C0(n5869), .Y(n1844)
         );
  OAI222XL U7891 ( .A0(n1834), .A1(n5719), .B0(n1835), .B1(n5691), .C0(n6482), 
        .C1(n5743), .Y(n1845) );
  OAI222XL U7892 ( .A0(n6400), .A1(n5875), .B0(n1800), .B1(n1787), .C0(n267), 
        .C1(n1788), .Y(n4165) );
  AOI211X1 U7893 ( .A0(n5925), .A1(n6483), .B0(n1801), .C0(n5869), .Y(n1800)
         );
  OAI222XL U7894 ( .A0(n1790), .A1(n5719), .B0(n1791), .B1(n5691), .C0(n6484), 
        .C1(n5743), .Y(n1801) );
  OAI222XL U7895 ( .A0(n6401), .A1(n5875), .B0(n1755), .B1(n1742), .C0(n259), 
        .C1(n1743), .Y(n4157) );
  AOI211X1 U7896 ( .A0(n5925), .A1(n6485), .B0(n1756), .C0(n5869), .Y(n1755)
         );
  OAI222XL U7897 ( .A0(n1745), .A1(n5720), .B0(n1746), .B1(n5691), .C0(n6486), 
        .C1(n5743), .Y(n1756) );
  OAI222XL U7898 ( .A0(n6402), .A1(n5875), .B0(n1711), .B1(n1698), .C0(n251), 
        .C1(n1699), .Y(n4149) );
  AOI211X1 U7899 ( .A0(n5925), .A1(n6487), .B0(n1712), .C0(n5869), .Y(n1711)
         );
  OAI222XL U7900 ( .A0(n1701), .A1(n5719), .B0(n1702), .B1(n5691), .C0(n6488), 
        .C1(n5743), .Y(n1712) );
  OAI222XL U7901 ( .A0(n6403), .A1(n5875), .B0(n1667), .B1(n1654), .C0(n243), 
        .C1(n1655), .Y(n4141) );
  AOI211X1 U7902 ( .A0(n5925), .A1(n6489), .B0(n1668), .C0(n5869), .Y(n1667)
         );
  OAI222XL U7903 ( .A0(n1657), .A1(n6501), .B0(n1658), .B1(n5691), .C0(n6490), 
        .C1(n5743), .Y(n1668) );
  OAI222XL U7904 ( .A0(n6404), .A1(n5875), .B0(n1623), .B1(n1610), .C0(n235), 
        .C1(n1611), .Y(n4133) );
  AOI211X1 U7905 ( .A0(n5925), .A1(n6491), .B0(n1624), .C0(n5869), .Y(n1623)
         );
  OAI222XL U7906 ( .A0(n1613), .A1(n5720), .B0(n1614), .B1(n5691), .C0(n6492), 
        .C1(n5743), .Y(n1624) );
  OAI222XL U7907 ( .A0(n6405), .A1(n5875), .B0(n1579), .B1(n1566), .C0(n227), 
        .C1(n1567), .Y(n4125) );
  AOI211X1 U7908 ( .A0(n5925), .A1(n6493), .B0(n1580), .C0(n5869), .Y(n1579)
         );
  OAI222XL U7909 ( .A0(n1569), .A1(n5718), .B0(n1570), .B1(n5691), .C0(n6494), 
        .C1(n5743), .Y(n1580) );
  OAI222XL U7910 ( .A0(n6406), .A1(n5872), .B0(n1535), .B1(n1522), .C0(n219), 
        .C1(n1523), .Y(n4117) );
  AOI211X1 U7911 ( .A0(n5925), .A1(n6495), .B0(n1536), .C0(n5869), .Y(n1535)
         );
  OAI222XL U7912 ( .A0(n1525), .A1(n5718), .B0(n1526), .B1(n5691), .C0(n6496), 
        .C1(n5743), .Y(n1536) );
  OAI222XL U7913 ( .A0(n6407), .A1(n5874), .B0(n1491), .B1(n1478), .C0(n211), 
        .C1(n1479), .Y(n4109) );
  OAI222XL U7914 ( .A0(n1481), .A1(n5718), .B0(n1482), .B1(n5693), .C0(n6498), 
        .C1(n5745), .Y(n1492) );
  OAI222XL U7915 ( .A0(n6347), .A1(n5883), .B0(n3941), .B1(n3929), .C0(n698), 
        .C1(n3930), .Y(n4596) );
  AOI211X1 U7916 ( .A0(n5929), .A1(n3931), .B0(n3942), .C0(n5876), .Y(n3941)
         );
  OAI222XL U7917 ( .A0(n3933), .A1(n5716), .B0(n3934), .B1(n5689), .C0(n6424), 
        .C1(n5742), .Y(n3942) );
  OAI222XL U7918 ( .A0(n6348), .A1(n5883), .B0(n3902), .B1(n3890), .C0(n690), 
        .C1(n3891), .Y(n4588) );
  AOI211X1 U7919 ( .A0(n5929), .A1(n3892), .B0(n3903), .C0(n5876), .Y(n3902)
         );
  OAI222XL U7920 ( .A0(n3894), .A1(n5716), .B0(n3895), .B1(n5690), .C0(n6425), 
        .C1(n5742), .Y(n3903) );
  OAI222XL U7921 ( .A0(n6349), .A1(n5883), .B0(n3863), .B1(n3851), .C0(n682), 
        .C1(n3852), .Y(n4580) );
  AOI211X1 U7922 ( .A0(n5929), .A1(n3853), .B0(n3864), .C0(n5876), .Y(n3863)
         );
  OAI222XL U7923 ( .A0(n3855), .A1(n5716), .B0(n3856), .B1(n5690), .C0(n6426), 
        .C1(n5742), .Y(n3864) );
  OAI222XL U7924 ( .A0(n6350), .A1(n5883), .B0(n3824), .B1(n3812), .C0(n674), 
        .C1(n3813), .Y(n4572) );
  AOI211X1 U7925 ( .A0(n5929), .A1(n3814), .B0(n3825), .C0(n5876), .Y(n3824)
         );
  OAI222XL U7926 ( .A0(n3816), .A1(n5717), .B0(n3817), .B1(n5690), .C0(n6427), 
        .C1(n5742), .Y(n3825) );
  OAI222XL U7927 ( .A0(n6351), .A1(n5883), .B0(n3785), .B1(n3773), .C0(n666), 
        .C1(n3774), .Y(n4564) );
  AOI211X1 U7928 ( .A0(n5929), .A1(n3775), .B0(n3786), .C0(n5876), .Y(n3785)
         );
  OAI222XL U7929 ( .A0(n3777), .A1(n5716), .B0(n3778), .B1(n5690), .C0(n6428), 
        .C1(n5742), .Y(n3786) );
  OAI222XL U7930 ( .A0(n6352), .A1(n5883), .B0(n3746), .B1(n3734), .C0(n658), 
        .C1(n3735), .Y(n4556) );
  AOI211X1 U7931 ( .A0(n5929), .A1(n3736), .B0(n3747), .C0(n5876), .Y(n3746)
         );
  OAI222XL U7932 ( .A0(n3738), .A1(n5717), .B0(n3739), .B1(n5689), .C0(n6429), 
        .C1(n5742), .Y(n3747) );
  OAI222XL U7933 ( .A0(n6353), .A1(n5883), .B0(n3702), .B1(n3690), .C0(n650), 
        .C1(n5670), .Y(n4548) );
  AOI211X1 U7934 ( .A0(n5929), .A1(n3692), .B0(n3703), .C0(n5876), .Y(n3702)
         );
  OAI222XL U7935 ( .A0(n3694), .A1(n5717), .B0(n3695), .B1(n6004), .C0(n6430), 
        .C1(n5742), .Y(n3703) );
  OAI222XL U7936 ( .A0(n6354), .A1(n5883), .B0(n3663), .B1(n3651), .C0(n642), 
        .C1(n3652), .Y(n4540) );
  AOI211X1 U7937 ( .A0(n5929), .A1(n3653), .B0(n3664), .C0(n5876), .Y(n3663)
         );
  OAI222XL U7938 ( .A0(n3655), .A1(n5716), .B0(n3656), .B1(n6067), .C0(n6431), 
        .C1(n5742), .Y(n3664) );
  OAI222XL U7939 ( .A0(n6355), .A1(n5883), .B0(n3624), .B1(n3612), .C0(n634), 
        .C1(n3613), .Y(n4532) );
  AOI211X1 U7940 ( .A0(n5929), .A1(n3614), .B0(n3625), .C0(n5876), .Y(n3624)
         );
  OAI222XL U7941 ( .A0(n3616), .A1(n5716), .B0(n3617), .B1(n5689), .C0(n6432), 
        .C1(n5742), .Y(n3625) );
  OAI222XL U7942 ( .A0(n6356), .A1(n5883), .B0(n3585), .B1(n3573), .C0(n626), 
        .C1(n3574), .Y(n4524) );
  AOI211X1 U7943 ( .A0(n5929), .A1(n3575), .B0(n3586), .C0(n5876), .Y(n3585)
         );
  OAI222XL U7944 ( .A0(n3577), .A1(n5717), .B0(n3578), .B1(n5689), .C0(n6433), 
        .C1(n5742), .Y(n3586) );
  OAI222XL U7945 ( .A0(n6357), .A1(n5883), .B0(n3546), .B1(n3534), .C0(n618), 
        .C1(n3535), .Y(n4516) );
  AOI211X1 U7946 ( .A0(n5929), .A1(n3536), .B0(n3547), .C0(n5876), .Y(n3546)
         );
  OAI222XL U7947 ( .A0(n3538), .A1(n5717), .B0(n3539), .B1(n5690), .C0(n6434), 
        .C1(n5742), .Y(n3547) );
  OAI222XL U7948 ( .A0(n6358), .A1(n5885), .B0(n3507), .B1(n3495), .C0(n610), 
        .C1(n3496), .Y(n4508) );
  AOI211X1 U7949 ( .A0(n5929), .A1(n3497), .B0(n3508), .C0(n5876), .Y(n3507)
         );
  OAI222XL U7950 ( .A0(n3499), .A1(n5715), .B0(n3500), .B1(n6420), .C0(n6435), 
        .C1(n5742), .Y(n3508) );
  OAI222XL U7951 ( .A0(n6359), .A1(n5884), .B0(n3468), .B1(n3456), .C0(n602), 
        .C1(n3457), .Y(n4500) );
  AOI211X1 U7952 ( .A0(n5929), .A1(n3458), .B0(n3469), .C0(n5877), .Y(n3468)
         );
  OAI222XL U7953 ( .A0(n3460), .A1(n5716), .B0(n3461), .B1(n6420), .C0(n6436), 
        .C1(n5742), .Y(n3469) );
  OAI222XL U7954 ( .A0(n6360), .A1(n5883), .B0(n3429), .B1(n3417), .C0(n594), 
        .C1(n3418), .Y(n4492) );
  AOI211X1 U7955 ( .A0(n5929), .A1(n3419), .B0(n3430), .C0(n5877), .Y(n3429)
         );
  OAI222XL U7956 ( .A0(n3421), .A1(n5715), .B0(n3422), .B1(n6420), .C0(n6437), 
        .C1(n5742), .Y(n3430) );
  OAI222XL U7957 ( .A0(n6361), .A1(n5885), .B0(n3385), .B1(n3373), .C0(n586), 
        .C1(n3374), .Y(n4484) );
  AOI211X1 U7958 ( .A0(n5929), .A1(n3375), .B0(n3386), .C0(n5877), .Y(n3385)
         );
  OAI222XL U7959 ( .A0(n3377), .A1(n5717), .B0(n3378), .B1(n6420), .C0(n6438), 
        .C1(n5742), .Y(n3386) );
  OAI222XL U7960 ( .A0(n6362), .A1(n5884), .B0(n3346), .B1(n3334), .C0(n578), 
        .C1(n3335), .Y(n4476) );
  AOI211X1 U7961 ( .A0(n5929), .A1(n3336), .B0(n3347), .C0(n5877), .Y(n3346)
         );
  OAI222XL U7962 ( .A0(n3338), .A1(n5717), .B0(n3339), .B1(n6420), .C0(n6439), 
        .C1(n5740), .Y(n3347) );
  OAI222XL U7963 ( .A0(n6363), .A1(n5883), .B0(n3307), .B1(n3295), .C0(n570), 
        .C1(n3296), .Y(n4468) );
  AOI211X1 U7964 ( .A0(n5929), .A1(n3297), .B0(n3308), .C0(n5877), .Y(n3307)
         );
  OAI222XL U7965 ( .A0(n3299), .A1(n5717), .B0(n3300), .B1(n6420), .C0(n6440), 
        .C1(n5742), .Y(n3308) );
  OAI222XL U7966 ( .A0(n6364), .A1(n5885), .B0(n3268), .B1(n3256), .C0(n562), 
        .C1(n3257), .Y(n4460) );
  AOI211X1 U7967 ( .A0(n5929), .A1(n3258), .B0(n3269), .C0(n5877), .Y(n3268)
         );
  OAI222XL U7968 ( .A0(n3260), .A1(n5715), .B0(n3261), .B1(n5690), .C0(n6441), 
        .C1(n5742), .Y(n3269) );
  OAI222XL U7969 ( .A0(n6365), .A1(n5884), .B0(n3229), .B1(n3217), .C0(n554), 
        .C1(n3218), .Y(n4452) );
  AOI211X1 U7970 ( .A0(n5929), .A1(n3219), .B0(n3230), .C0(n5877), .Y(n3229)
         );
  OAI222XL U7971 ( .A0(n3221), .A1(n5715), .B0(n3222), .B1(n5690), .C0(n6442), 
        .C1(n5741), .Y(n3230) );
  OAI222XL U7972 ( .A0(n6366), .A1(n5883), .B0(n3190), .B1(n3178), .C0(n546), 
        .C1(n3179), .Y(n4444) );
  AOI211X1 U7973 ( .A0(n5929), .A1(n3180), .B0(n3191), .C0(n5877), .Y(n3190)
         );
  OAI222XL U7974 ( .A0(n3182), .A1(n5717), .B0(n3183), .B1(n5690), .C0(n6443), 
        .C1(n5740), .Y(n3191) );
  OAI222XL U7975 ( .A0(n6367), .A1(n5883), .B0(n3151), .B1(n3139), .C0(n538), 
        .C1(n4674), .Y(n4436) );
  AOI211X1 U7976 ( .A0(n5929), .A1(n3141), .B0(n3152), .C0(n5877), .Y(n3151)
         );
  OAI222XL U7977 ( .A0(n3143), .A1(n5715), .B0(n3144), .B1(n5690), .C0(n6444), 
        .C1(n5742), .Y(n3152) );
  OAI222XL U7978 ( .A0(n6368), .A1(n5885), .B0(n3112), .B1(n3100), .C0(n530), 
        .C1(n3101), .Y(n4428) );
  AOI211X1 U7979 ( .A0(n5929), .A1(n3102), .B0(n3113), .C0(n5877), .Y(n3112)
         );
  OAI222XL U7980 ( .A0(n3104), .A1(n5715), .B0(n3105), .B1(n5690), .C0(n6445), 
        .C1(n5740), .Y(n3113) );
  OAI222XL U7981 ( .A0(n6369), .A1(n5884), .B0(n3068), .B1(n3056), .C0(n522), 
        .C1(n3057), .Y(n4420) );
  AOI211X1 U7982 ( .A0(n5929), .A1(n3058), .B0(n3069), .C0(n5877), .Y(n3068)
         );
  OAI222XL U7983 ( .A0(n3060), .A1(n5715), .B0(n3061), .B1(n5690), .C0(n6446), 
        .C1(n5741), .Y(n3069) );
  OAI222XL U7984 ( .A0(n6370), .A1(n5884), .B0(n3029), .B1(n3017), .C0(n514), 
        .C1(n3018), .Y(n4412) );
  AOI211X1 U7985 ( .A0(n5929), .A1(n3019), .B0(n3030), .C0(n5877), .Y(n3029)
         );
  OAI222XL U7986 ( .A0(n3021), .A1(n5715), .B0(n3022), .B1(n5690), .C0(n6447), 
        .C1(n5740), .Y(n3030) );
  OAI222XL U7987 ( .A0(n6371), .A1(n5884), .B0(n2990), .B1(n2978), .C0(n506), 
        .C1(n2979), .Y(n4404) );
  AOI211X1 U7988 ( .A0(n5929), .A1(n2980), .B0(n2991), .C0(n5877), .Y(n2990)
         );
  OAI222XL U7989 ( .A0(n2982), .A1(n5715), .B0(n2983), .B1(n5690), .C0(n6448), 
        .C1(n5740), .Y(n2991) );
  OAI222XL U7990 ( .A0(n6372), .A1(n5884), .B0(n2951), .B1(n2939), .C0(n498), 
        .C1(n4675), .Y(n4396) );
  AOI211X1 U7991 ( .A0(n5929), .A1(n2941), .B0(n2952), .C0(n5878), .Y(n2951)
         );
  OAI222XL U7992 ( .A0(n2943), .A1(n5715), .B0(n2944), .B1(n5690), .C0(n6449), 
        .C1(n5742), .Y(n2952) );
  OAI222XL U7993 ( .A0(n6373), .A1(n5884), .B0(n2912), .B1(n2900), .C0(n490), 
        .C1(n2901), .Y(n4388) );
  AOI211X1 U7994 ( .A0(n5929), .A1(n2902), .B0(n2913), .C0(n5878), .Y(n2912)
         );
  OAI222XL U7995 ( .A0(n2904), .A1(n5715), .B0(n2905), .B1(n5690), .C0(n6450), 
        .C1(n5740), .Y(n2913) );
  OAI222XL U7996 ( .A0(n6374), .A1(n5884), .B0(n2873), .B1(n2861), .C0(n482), 
        .C1(n2862), .Y(n4380) );
  AOI211X1 U7997 ( .A0(n5929), .A1(n2863), .B0(n2874), .C0(n5878), .Y(n2873)
         );
  OAI222XL U7998 ( .A0(n2865), .A1(n5715), .B0(n2866), .B1(n5690), .C0(n6451), 
        .C1(n5740), .Y(n2874) );
  OAI222XL U7999 ( .A0(n6375), .A1(n5884), .B0(n2834), .B1(n2822), .C0(n474), 
        .C1(n2823), .Y(n4372) );
  AOI211X1 U8000 ( .A0(n5929), .A1(n2824), .B0(n2835), .C0(n5878), .Y(n2834)
         );
  OAI222XL U8001 ( .A0(n2826), .A1(n5715), .B0(n2827), .B1(n5690), .C0(n6452), 
        .C1(n5740), .Y(n2835) );
  OAI222XL U8002 ( .A0(n6376), .A1(n5884), .B0(n2795), .B1(n2783), .C0(n466), 
        .C1(n2784), .Y(n4364) );
  AOI211X1 U8003 ( .A0(n5928), .A1(n2785), .B0(n2796), .C0(n5878), .Y(n2795)
         );
  OAI222XL U8004 ( .A0(n2787), .A1(n5715), .B0(n2788), .B1(n5690), .C0(n6453), 
        .C1(n5742), .Y(n2796) );
  OAI222XL U8005 ( .A0(n6377), .A1(n5884), .B0(n2751), .B1(n2739), .C0(n458), 
        .C1(n2740), .Y(n4356) );
  AOI211X1 U8006 ( .A0(n5928), .A1(n2741), .B0(n2752), .C0(n5878), .Y(n2751)
         );
  OAI222XL U8007 ( .A0(n2743), .A1(n5715), .B0(n2744), .B1(n5690), .C0(n6454), 
        .C1(n5742), .Y(n2752) );
  OAI222XL U8008 ( .A0(n6378), .A1(n5884), .B0(n2712), .B1(n2700), .C0(n450), 
        .C1(n2701), .Y(n4348) );
  AOI211X1 U8009 ( .A0(n5928), .A1(n2702), .B0(n2713), .C0(n5878), .Y(n2712)
         );
  OAI222XL U8010 ( .A0(n2704), .A1(n5715), .B0(n2705), .B1(n5690), .C0(n6455), 
        .C1(n5742), .Y(n2713) );
  OAI222XL U8011 ( .A0(n6379), .A1(n5884), .B0(n2673), .B1(n2661), .C0(n442), 
        .C1(n2662), .Y(n4340) );
  AOI211X1 U8012 ( .A0(n5928), .A1(n2663), .B0(n2674), .C0(n5878), .Y(n2673)
         );
  OAI222XL U8013 ( .A0(n2665), .A1(n5715), .B0(n2666), .B1(n5689), .C0(n6456), 
        .C1(n5742), .Y(n2674) );
  OAI222XL U8014 ( .A0(n6380), .A1(n5884), .B0(n2634), .B1(n2622), .C0(n434), 
        .C1(n2623), .Y(n4332) );
  AOI211X1 U8015 ( .A0(n5928), .A1(n2624), .B0(n2635), .C0(n5878), .Y(n2634)
         );
  OAI222XL U8016 ( .A0(n2626), .A1(n5715), .B0(n2627), .B1(n5689), .C0(n6457), 
        .C1(n5742), .Y(n2635) );
  OAI222XL U8017 ( .A0(n6381), .A1(n5884), .B0(n2595), .B1(n2583), .C0(n426), 
        .C1(n2584), .Y(n4324) );
  AOI211X1 U8018 ( .A0(n5928), .A1(n2585), .B0(n2596), .C0(n5878), .Y(n2595)
         );
  OAI222XL U8019 ( .A0(n2587), .A1(n5715), .B0(n2588), .B1(n5689), .C0(n6458), 
        .C1(n5742), .Y(n2596) );
  OAI222XL U8020 ( .A0(n6382), .A1(n5885), .B0(n2556), .B1(n2544), .C0(n418), 
        .C1(n2545), .Y(n4316) );
  AOI211X1 U8021 ( .A0(n5928), .A1(n2546), .B0(n2557), .C0(n5878), .Y(n2556)
         );
  OAI222XL U8022 ( .A0(n2548), .A1(n5716), .B0(n2549), .B1(n5689), .C0(n6459), 
        .C1(n5742), .Y(n2557) );
  OAI222XL U8023 ( .A0(n6383), .A1(n5885), .B0(n2517), .B1(n2505), .C0(n410), 
        .C1(n2506), .Y(n4308) );
  AOI211X1 U8024 ( .A0(n5928), .A1(n2507), .B0(n2518), .C0(n5878), .Y(n2517)
         );
  OAI222XL U8025 ( .A0(n2509), .A1(n5716), .B0(n2510), .B1(n5689), .C0(n6460), 
        .C1(n5742), .Y(n2518) );
  OAI222XL U8026 ( .A0(n6384), .A1(n5885), .B0(n2478), .B1(n2466), .C0(n402), 
        .C1(n2467), .Y(n4300) );
  AOI211X1 U8027 ( .A0(n5928), .A1(n2468), .B0(n2479), .C0(n5878), .Y(n2478)
         );
  OAI222XL U8028 ( .A0(n2470), .A1(n5716), .B0(n2471), .B1(n5689), .C0(n6461), 
        .C1(n5742), .Y(n2479) );
  OAI222XL U8029 ( .A0(n6385), .A1(n5885), .B0(n2434), .B1(n2422), .C0(n394), 
        .C1(n2423), .Y(n4292) );
  AOI211X1 U8030 ( .A0(n5928), .A1(n2424), .B0(n2435), .C0(n5879), .Y(n2434)
         );
  OAI222XL U8031 ( .A0(n2426), .A1(n5716), .B0(n2427), .B1(n5689), .C0(n6462), 
        .C1(n5742), .Y(n2435) );
  OAI222XL U8032 ( .A0(n6386), .A1(n5885), .B0(n2395), .B1(n2383), .C0(n386), 
        .C1(n2384), .Y(n4284) );
  AOI211X1 U8033 ( .A0(n5928), .A1(n2385), .B0(n2396), .C0(n5879), .Y(n2395)
         );
  OAI222XL U8034 ( .A0(n2387), .A1(n5716), .B0(n2388), .B1(n5689), .C0(n6463), 
        .C1(n5742), .Y(n2396) );
  OAI222XL U8035 ( .A0(n6387), .A1(n5885), .B0(n2356), .B1(n2344), .C0(n378), 
        .C1(n2345), .Y(n4276) );
  AOI211X1 U8036 ( .A0(n5928), .A1(n2346), .B0(n2357), .C0(n5876), .Y(n2356)
         );
  OAI222XL U8037 ( .A0(n2348), .A1(n5716), .B0(n2349), .B1(n5689), .C0(n6464), 
        .C1(n5742), .Y(n2357) );
  OAI222XL U8038 ( .A0(n6388), .A1(n5885), .B0(n2317), .B1(n2305), .C0(n370), 
        .C1(n2306), .Y(n4268) );
  AOI211X1 U8039 ( .A0(n5928), .A1(n2307), .B0(n2318), .C0(n5879), .Y(n2317)
         );
  OAI222XL U8040 ( .A0(n2309), .A1(n5716), .B0(n2310), .B1(n5689), .C0(n6465), 
        .C1(n5742), .Y(n2318) );
  OAI222XL U8041 ( .A0(n6389), .A1(n5885), .B0(n2278), .B1(n2266), .C0(n362), 
        .C1(n2267), .Y(n4260) );
  AOI211X1 U8042 ( .A0(n5928), .A1(n2268), .B0(n2279), .C0(n5876), .Y(n2278)
         );
  OAI222XL U8043 ( .A0(n2270), .A1(n5716), .B0(n2271), .B1(n5689), .C0(n6466), 
        .C1(n5742), .Y(n2279) );
  OAI222XL U8044 ( .A0(n6390), .A1(n5885), .B0(n2239), .B1(n2227), .C0(n354), 
        .C1(n2228), .Y(n4252) );
  AOI211X1 U8045 ( .A0(n5928), .A1(n2229), .B0(n2240), .C0(n5879), .Y(n2239)
         );
  OAI222XL U8046 ( .A0(n2231), .A1(n5716), .B0(n2232), .B1(n5689), .C0(n6467), 
        .C1(n5742), .Y(n2240) );
  OAI222XL U8047 ( .A0(n6391), .A1(n5885), .B0(n2200), .B1(n2188), .C0(n346), 
        .C1(n2189), .Y(n4244) );
  AOI211X1 U8048 ( .A0(n5928), .A1(n2190), .B0(n2201), .C0(n5876), .Y(n2200)
         );
  OAI222XL U8049 ( .A0(n2192), .A1(n5716), .B0(n2193), .B1(n5689), .C0(n6468), 
        .C1(n5742), .Y(n2201) );
  OAI222XL U8050 ( .A0(n6392), .A1(n5885), .B0(n2161), .B1(n2149), .C0(n338), 
        .C1(n2150), .Y(n4236) );
  AOI211X1 U8051 ( .A0(n5928), .A1(n2151), .B0(n2162), .C0(n5879), .Y(n2161)
         );
  OAI222XL U8052 ( .A0(n2153), .A1(n5716), .B0(n2154), .B1(n5689), .C0(n6469), 
        .C1(n5742), .Y(n2162) );
  OAI222XL U8053 ( .A0(n6393), .A1(n5885), .B0(n2117), .B1(n2105), .C0(n330), 
        .C1(n2106), .Y(n4228) );
  AOI211X1 U8054 ( .A0(n5928), .A1(n2107), .B0(n2118), .C0(n5876), .Y(n2117)
         );
  OAI222XL U8055 ( .A0(n2109), .A1(n5716), .B0(n2110), .B1(n5689), .C0(n6470), 
        .C1(n5742), .Y(n2118) );
  OAI222XL U8056 ( .A0(n6394), .A1(n5883), .B0(n2078), .B1(n2066), .C0(n322), 
        .C1(n2067), .Y(n4220) );
  AOI211X1 U8057 ( .A0(n5928), .A1(n2068), .B0(n2079), .C0(n5876), .Y(n2078)
         );
  OAI222XL U8058 ( .A0(n2070), .A1(n5717), .B0(n2071), .B1(n5689), .C0(n6471), 
        .C1(n5742), .Y(n2079) );
  OAI222XL U8059 ( .A0(n6395), .A1(n5883), .B0(n2039), .B1(n2027), .C0(n314), 
        .C1(n2028), .Y(n4212) );
  AOI211X1 U8060 ( .A0(n5928), .A1(n2029), .B0(n2040), .C0(n5879), .Y(n2039)
         );
  OAI222XL U8061 ( .A0(n2031), .A1(n5717), .B0(n2032), .B1(n5688), .C0(n6472), 
        .C1(n5742), .Y(n2040) );
  OAI222XL U8062 ( .A0(n6396), .A1(n5885), .B0(n1998), .B1(n1987), .C0(n306), 
        .C1(n1988), .Y(n4204) );
  AOI211X1 U8063 ( .A0(n5928), .A1(n6473), .B0(n1999), .C0(n5879), .Y(n1998)
         );
  OAI222XL U8064 ( .A0(n1990), .A1(n5717), .B0(n1991), .B1(n5688), .C0(n6474), 
        .C1(n5741), .Y(n1999) );
  OAI222XL U8065 ( .A0(n6397), .A1(n5885), .B0(n1959), .B1(n1948), .C0(n298), 
        .C1(n1949), .Y(n4196) );
  AOI211X1 U8066 ( .A0(n5928), .A1(n6475), .B0(n1960), .C0(n5876), .Y(n1959)
         );
  OAI222XL U8067 ( .A0(n1951), .A1(n5717), .B0(n1952), .B1(n5688), .C0(n6476), 
        .C1(n5740), .Y(n1960) );
  OAI222XL U8068 ( .A0(n6398), .A1(n5885), .B0(n1920), .B1(n1909), .C0(n290), 
        .C1(n1910), .Y(n4188) );
  AOI211X1 U8069 ( .A0(n5928), .A1(n6477), .B0(n1921), .C0(n5879), .Y(n1920)
         );
  OAI222XL U8070 ( .A0(n1912), .A1(n5717), .B0(n1913), .B1(n5688), .C0(n6478), 
        .C1(n5740), .Y(n1921) );
  OAI222XL U8071 ( .A0(n4832), .A1(n5884), .B0(n1881), .B1(n1870), .C0(n282), 
        .C1(n1871), .Y(n4180) );
  AOI211X1 U8072 ( .A0(n5928), .A1(n6479), .B0(n1882), .C0(n5879), .Y(n1881)
         );
  OAI222XL U8073 ( .A0(n1873), .A1(n5717), .B0(n1874), .B1(n5688), .C0(n6480), 
        .C1(n5740), .Y(n1882) );
  OAI222XL U8074 ( .A0(n6399), .A1(n5884), .B0(n1842), .B1(n1831), .C0(n274), 
        .C1(n4643), .Y(n4172) );
  AOI211X1 U8075 ( .A0(n5928), .A1(n6481), .B0(n1843), .C0(n5879), .Y(n1842)
         );
  OAI222XL U8076 ( .A0(n1834), .A1(n5717), .B0(n1835), .B1(n5688), .C0(n6482), 
        .C1(n5740), .Y(n1843) );
  OAI222XL U8077 ( .A0(n6400), .A1(n5884), .B0(n1798), .B1(n1787), .C0(n266), 
        .C1(n1788), .Y(n4164) );
  AOI211X1 U8078 ( .A0(n5928), .A1(n6483), .B0(n1799), .C0(n5879), .Y(n1798)
         );
  OAI222XL U8079 ( .A0(n1790), .A1(n5717), .B0(n1791), .B1(n5688), .C0(n6484), 
        .C1(n5741), .Y(n1799) );
  OAI222XL U8080 ( .A0(n6401), .A1(n5883), .B0(n1753), .B1(n1742), .C0(n258), 
        .C1(n1743), .Y(n4156) );
  AOI211X1 U8081 ( .A0(n5928), .A1(n6485), .B0(n1754), .C0(n5879), .Y(n1753)
         );
  OAI222XL U8082 ( .A0(n1745), .A1(n5717), .B0(n1746), .B1(n5688), .C0(n6486), 
        .C1(n5740), .Y(n1754) );
  OAI222XL U8083 ( .A0(n6402), .A1(n5885), .B0(n1709), .B1(n1698), .C0(n250), 
        .C1(n1699), .Y(n4148) );
  AOI211X1 U8084 ( .A0(n5928), .A1(n6487), .B0(n1710), .C0(n5879), .Y(n1709)
         );
  OAI222XL U8085 ( .A0(n1701), .A1(n5717), .B0(n1702), .B1(n5688), .C0(n6488), 
        .C1(n5740), .Y(n1710) );
  OAI222XL U8086 ( .A0(n6403), .A1(n5884), .B0(n1665), .B1(n1654), .C0(n242), 
        .C1(n1655), .Y(n4140) );
  AOI211X1 U8087 ( .A0(n5928), .A1(n6489), .B0(n1666), .C0(n5879), .Y(n1665)
         );
  OAI222XL U8088 ( .A0(n1657), .A1(n5717), .B0(n1658), .B1(n5688), .C0(n6490), 
        .C1(n5741), .Y(n1666) );
  OAI222XL U8089 ( .A0(n6404), .A1(n5884), .B0(n1621), .B1(n1610), .C0(n234), 
        .C1(n1611), .Y(n4132) );
  AOI211X1 U8090 ( .A0(n5928), .A1(n6491), .B0(n1622), .C0(n5879), .Y(n1621)
         );
  OAI222XL U8091 ( .A0(n1613), .A1(n5717), .B0(n1614), .B1(n5688), .C0(n6492), 
        .C1(n5740), .Y(n1622) );
  OAI222XL U8092 ( .A0(n6405), .A1(n5883), .B0(n1577), .B1(n1566), .C0(n226), 
        .C1(n1567), .Y(n4124) );
  AOI211X1 U8093 ( .A0(n5928), .A1(n6493), .B0(n1578), .C0(n5879), .Y(n1577)
         );
  OAI222XL U8094 ( .A0(n1569), .A1(n5716), .B0(n1570), .B1(n5688), .C0(n6494), 
        .C1(n5740), .Y(n1578) );
  OAI222XL U8095 ( .A0(n6406), .A1(n5883), .B0(n1533), .B1(n1522), .C0(n218), 
        .C1(n1523), .Y(n4116) );
  AOI211X1 U8096 ( .A0(n5928), .A1(n6495), .B0(n1534), .C0(n5879), .Y(n1533)
         );
  OAI222XL U8097 ( .A0(n1525), .A1(n5715), .B0(n1526), .B1(n5688), .C0(n6496), 
        .C1(n5741), .Y(n1534) );
  OAI222XL U8098 ( .A0(n6407), .A1(n5885), .B0(n1489), .B1(n1478), .C0(n210), 
        .C1(n1479), .Y(n4108) );
  OAI222XL U8099 ( .A0(n1481), .A1(n5715), .B0(n1482), .B1(n5690), .C0(n6498), 
        .C1(n5742), .Y(n1490) );
  OAI222XL U8100 ( .A0(n3933), .A1(n5711), .B0(n3934), .B1(n5685), .C0(n6424), 
        .C1(n5738), .Y(n3940) );
  OAI222XL U8101 ( .A0(n6348), .A1(n5894), .B0(n3900), .B1(n3890), .C0(n689), 
        .C1(n3891), .Y(n4587) );
  AOI211X1 U8102 ( .A0(n5935), .A1(n3892), .B0(n3901), .C0(n5889), .Y(n3900)
         );
  OAI222XL U8103 ( .A0(n3894), .A1(n5713), .B0(n3895), .B1(n5687), .C0(n6425), 
        .C1(n5738), .Y(n3901) );
  OAI222XL U8104 ( .A0(n6349), .A1(n5895), .B0(n3861), .B1(n3851), .C0(n681), 
        .C1(n3852), .Y(n4579) );
  AOI211X1 U8105 ( .A0(n5935), .A1(n3853), .B0(n3862), .C0(n5889), .Y(n3861)
         );
  OAI222XL U8106 ( .A0(n3855), .A1(n5713), .B0(n3856), .B1(n5687), .C0(n6426), 
        .C1(n5739), .Y(n3862) );
  OAI222XL U8107 ( .A0(n6350), .A1(n5893), .B0(n3822), .B1(n3812), .C0(n673), 
        .C1(n3813), .Y(n4571) );
  AOI211X1 U8108 ( .A0(n5935), .A1(n3814), .B0(n3823), .C0(n5889), .Y(n3822)
         );
  OAI222XL U8109 ( .A0(n3816), .A1(n5714), .B0(n3817), .B1(n5687), .C0(n6427), 
        .C1(n5739), .Y(n3823) );
  OAI222XL U8110 ( .A0(n6351), .A1(n5894), .B0(n3783), .B1(n3773), .C0(n665), 
        .C1(n3774), .Y(n4563) );
  AOI211X1 U8111 ( .A0(n5935), .A1(n3775), .B0(n3784), .C0(n5889), .Y(n3783)
         );
  OAI222XL U8112 ( .A0(n3777), .A1(n5712), .B0(n3778), .B1(n5687), .C0(n6428), 
        .C1(n5739), .Y(n3784) );
  OAI222XL U8113 ( .A0(n6352), .A1(n5895), .B0(n3744), .B1(n3734), .C0(n657), 
        .C1(n3735), .Y(n4555) );
  AOI211X1 U8114 ( .A0(n5935), .A1(n3736), .B0(n3745), .C0(n5889), .Y(n3744)
         );
  OAI222XL U8115 ( .A0(n3738), .A1(n5712), .B0(n3739), .B1(n5687), .C0(n6429), 
        .C1(n5739), .Y(n3745) );
  OAI222XL U8116 ( .A0(n6353), .A1(n5893), .B0(n3700), .B1(n3690), .C0(n649), 
        .C1(n5670), .Y(n4547) );
  AOI211X1 U8117 ( .A0(n5935), .A1(n3692), .B0(n3701), .C0(n5889), .Y(n3700)
         );
  OAI222XL U8118 ( .A0(n3694), .A1(n5711), .B0(n3695), .B1(n5687), .C0(n6430), 
        .C1(n5739), .Y(n3701) );
  OAI222XL U8119 ( .A0(n6354), .A1(n5894), .B0(n3661), .B1(n3651), .C0(n641), 
        .C1(n3652), .Y(n4539) );
  AOI211X1 U8120 ( .A0(n5935), .A1(n3653), .B0(n3662), .C0(n5889), .Y(n3661)
         );
  OAI222XL U8121 ( .A0(n3655), .A1(n5711), .B0(n3656), .B1(n5687), .C0(n6431), 
        .C1(n5739), .Y(n3662) );
  OAI222XL U8122 ( .A0(n6355), .A1(n5895), .B0(n3622), .B1(n3612), .C0(n633), 
        .C1(n3613), .Y(n4531) );
  AOI211X1 U8123 ( .A0(n5935), .A1(n3614), .B0(n3623), .C0(n5889), .Y(n3622)
         );
  OAI222XL U8124 ( .A0(n3616), .A1(n5711), .B0(n3617), .B1(n5687), .C0(n6432), 
        .C1(n5739), .Y(n3623) );
  OAI222XL U8125 ( .A0(n6356), .A1(n5893), .B0(n3583), .B1(n3573), .C0(n625), 
        .C1(n3574), .Y(n4523) );
  AOI211X1 U8126 ( .A0(n5935), .A1(n3575), .B0(n3584), .C0(n5889), .Y(n3583)
         );
  OAI222XL U8127 ( .A0(n3577), .A1(n5711), .B0(n3578), .B1(n5687), .C0(n6433), 
        .C1(n5739), .Y(n3584) );
  OAI222XL U8128 ( .A0(n6357), .A1(n5894), .B0(n3544), .B1(n3534), .C0(n617), 
        .C1(n3535), .Y(n4515) );
  AOI211X1 U8129 ( .A0(n5935), .A1(n3536), .B0(n3545), .C0(n5889), .Y(n3544)
         );
  OAI222XL U8130 ( .A0(n3538), .A1(n5711), .B0(n3539), .B1(n5687), .C0(n6434), 
        .C1(n5739), .Y(n3545) );
  OAI222XL U8131 ( .A0(n6358), .A1(n5893), .B0(n3505), .B1(n3495), .C0(n609), 
        .C1(n3496), .Y(n4507) );
  AOI211X1 U8132 ( .A0(n5935), .A1(n3497), .B0(n3506), .C0(n5889), .Y(n3505)
         );
  OAI222XL U8133 ( .A0(n3499), .A1(n5712), .B0(n3500), .B1(n5687), .C0(n6435), 
        .C1(n5739), .Y(n3506) );
  OAI222XL U8134 ( .A0(n6359), .A1(n5893), .B0(n3466), .B1(n3456), .C0(n601), 
        .C1(n3457), .Y(n4499) );
  AOI211X1 U8135 ( .A0(n5935), .A1(n3458), .B0(n3467), .C0(n5886), .Y(n3466)
         );
  OAI222XL U8136 ( .A0(n3460), .A1(n5712), .B0(n3461), .B1(n5687), .C0(n6436), 
        .C1(n5739), .Y(n3467) );
  OAI222XL U8137 ( .A0(n6360), .A1(n5893), .B0(n3427), .B1(n3417), .C0(n593), 
        .C1(n3418), .Y(n4491) );
  AOI211X1 U8138 ( .A0(n5935), .A1(n3419), .B0(n3428), .C0(n5886), .Y(n3427)
         );
  OAI222XL U8139 ( .A0(n3421), .A1(n5712), .B0(n3422), .B1(n5687), .C0(n6437), 
        .C1(n5739), .Y(n3428) );
  OAI222XL U8140 ( .A0(n6361), .A1(n5893), .B0(n3383), .B1(n3373), .C0(n585), 
        .C1(n3374), .Y(n4483) );
  AOI211X1 U8141 ( .A0(n5935), .A1(n3375), .B0(n3384), .C0(n5886), .Y(n3383)
         );
  OAI222XL U8142 ( .A0(n3377), .A1(n5712), .B0(n3378), .B1(n5687), .C0(n6438), 
        .C1(n5739), .Y(n3384) );
  OAI222XL U8143 ( .A0(n6362), .A1(n5893), .B0(n3344), .B1(n3334), .C0(n577), 
        .C1(n3335), .Y(n4475) );
  AOI211X1 U8144 ( .A0(n5935), .A1(n3336), .B0(n3345), .C0(n5886), .Y(n3344)
         );
  OAI222XL U8145 ( .A0(n3338), .A1(n5712), .B0(n3339), .B1(n5687), .C0(n6439), 
        .C1(n5739), .Y(n3345) );
  OAI222XL U8146 ( .A0(n6363), .A1(n5893), .B0(n3305), .B1(n3295), .C0(n569), 
        .C1(n3296), .Y(n4467) );
  AOI211X1 U8147 ( .A0(n5935), .A1(n3297), .B0(n3306), .C0(n5886), .Y(n3305)
         );
  OAI222XL U8148 ( .A0(n3299), .A1(n5712), .B0(n3300), .B1(n5687), .C0(n6440), 
        .C1(n5739), .Y(n3306) );
  OAI222XL U8149 ( .A0(n6364), .A1(n5893), .B0(n3266), .B1(n3256), .C0(n561), 
        .C1(n3257), .Y(n4459) );
  AOI211X1 U8150 ( .A0(n5935), .A1(n3258), .B0(n3267), .C0(n5886), .Y(n3266)
         );
  OAI222XL U8151 ( .A0(n3260), .A1(n5712), .B0(n3261), .B1(n5686), .C0(n6441), 
        .C1(n5739), .Y(n3267) );
  OAI222XL U8152 ( .A0(n6365), .A1(n5893), .B0(n3227), .B1(n3217), .C0(n553), 
        .C1(n3218), .Y(n4451) );
  AOI211X1 U8153 ( .A0(n5935), .A1(n3219), .B0(n3228), .C0(n5886), .Y(n3227)
         );
  OAI222XL U8154 ( .A0(n3221), .A1(n5712), .B0(n3222), .B1(n5686), .C0(n6442), 
        .C1(n5739), .Y(n3228) );
  OAI222XL U8155 ( .A0(n6366), .A1(n5893), .B0(n3188), .B1(n3178), .C0(n545), 
        .C1(n3179), .Y(n4443) );
  AOI211X1 U8156 ( .A0(n5935), .A1(n3180), .B0(n3189), .C0(n5886), .Y(n3188)
         );
  OAI222XL U8157 ( .A0(n3182), .A1(n5712), .B0(n3183), .B1(n5686), .C0(n6443), 
        .C1(n5739), .Y(n3189) );
  OAI222XL U8158 ( .A0(n3143), .A1(n5712), .B0(n3144), .B1(n5686), .C0(n6444), 
        .C1(n5739), .Y(n3150) );
  OAI222XL U8159 ( .A0(n6368), .A1(n5893), .B0(n3110), .B1(n3100), .C0(n529), 
        .C1(n3101), .Y(n4427) );
  AOI211X1 U8160 ( .A0(n5935), .A1(n3102), .B0(n3111), .C0(n5886), .Y(n3110)
         );
  OAI222XL U8161 ( .A0(n3104), .A1(n5712), .B0(n3105), .B1(n5686), .C0(n6445), 
        .C1(n5739), .Y(n3111) );
  OAI222XL U8162 ( .A0(n6369), .A1(n5893), .B0(n3066), .B1(n3056), .C0(n521), 
        .C1(n3057), .Y(n4419) );
  AOI211X1 U8163 ( .A0(n5935), .A1(n3058), .B0(n3067), .C0(n5886), .Y(n3066)
         );
  OAI222XL U8164 ( .A0(n3060), .A1(n5712), .B0(n3061), .B1(n5686), .C0(n6446), 
        .C1(n5739), .Y(n3067) );
  OAI222XL U8165 ( .A0(n6370), .A1(n5894), .B0(n3027), .B1(n3017), .C0(n513), 
        .C1(n3018), .Y(n4411) );
  AOI211X1 U8166 ( .A0(n5935), .A1(n3019), .B0(n3028), .C0(n5886), .Y(n3027)
         );
  OAI222XL U8167 ( .A0(n3021), .A1(n5713), .B0(n3022), .B1(n5686), .C0(n6447), 
        .C1(n5737), .Y(n3028) );
  OAI222XL U8168 ( .A0(n6371), .A1(n5894), .B0(n2988), .B1(n2978), .C0(n505), 
        .C1(n2979), .Y(n4403) );
  AOI211X1 U8169 ( .A0(n5935), .A1(n2980), .B0(n2989), .C0(n5886), .Y(n2988)
         );
  OAI222XL U8170 ( .A0(n2982), .A1(n5713), .B0(n2983), .B1(n5686), .C0(n6448), 
        .C1(n5737), .Y(n2989) );
  OAI222XL U8171 ( .A0(n2943), .A1(n5713), .B0(n2944), .B1(n5686), .C0(n6449), 
        .C1(n5738), .Y(n2950) );
  OAI222XL U8172 ( .A0(n6373), .A1(n5894), .B0(n2910), .B1(n2900), .C0(n489), 
        .C1(n2901), .Y(n4387) );
  AOI211X1 U8173 ( .A0(n5935), .A1(n2902), .B0(n2911), .C0(n5887), .Y(n2910)
         );
  OAI222XL U8174 ( .A0(n2904), .A1(n5713), .B0(n2905), .B1(n5686), .C0(n6450), 
        .C1(n5737), .Y(n2911) );
  OAI222XL U8175 ( .A0(n6374), .A1(n5894), .B0(n2871), .B1(n2861), .C0(n481), 
        .C1(n2862), .Y(n4379) );
  AOI211X1 U8176 ( .A0(n5935), .A1(n2863), .B0(n2872), .C0(n5887), .Y(n2871)
         );
  OAI222XL U8177 ( .A0(n2865), .A1(n5713), .B0(n2866), .B1(n5686), .C0(n6451), 
        .C1(n6506), .Y(n2872) );
  OAI222XL U8178 ( .A0(n6375), .A1(n5894), .B0(n2832), .B1(n2822), .C0(n473), 
        .C1(n2823), .Y(n4371) );
  AOI211X1 U8179 ( .A0(n5935), .A1(n2824), .B0(n2833), .C0(n5887), .Y(n2832)
         );
  OAI222XL U8180 ( .A0(n2826), .A1(n5713), .B0(n2827), .B1(n5686), .C0(n6452), 
        .C1(n6506), .Y(n2833) );
  OAI222XL U8181 ( .A0(n6376), .A1(n5894), .B0(n2793), .B1(n2783), .C0(n465), 
        .C1(n2784), .Y(n4363) );
  AOI211X1 U8182 ( .A0(n5934), .A1(n2785), .B0(n2794), .C0(n5887), .Y(n2793)
         );
  OAI222XL U8183 ( .A0(n2787), .A1(n5713), .B0(n2788), .B1(n5686), .C0(n6453), 
        .C1(n6506), .Y(n2794) );
  OAI222XL U8184 ( .A0(n6377), .A1(n5894), .B0(n2749), .B1(n2739), .C0(n457), 
        .C1(n2740), .Y(n4355) );
  AOI211X1 U8185 ( .A0(n5934), .A1(n2741), .B0(n2750), .C0(n5887), .Y(n2749)
         );
  OAI222XL U8186 ( .A0(n2743), .A1(n5713), .B0(n2744), .B1(n5686), .C0(n6454), 
        .C1(n6506), .Y(n2750) );
  OAI222XL U8187 ( .A0(n6378), .A1(n5894), .B0(n2710), .B1(n2700), .C0(n449), 
        .C1(n2701), .Y(n4347) );
  AOI211X1 U8188 ( .A0(n5934), .A1(n2702), .B0(n2711), .C0(n5887), .Y(n2710)
         );
  OAI222XL U8189 ( .A0(n2704), .A1(n5713), .B0(n2705), .B1(n5686), .C0(n6455), 
        .C1(n6506), .Y(n2711) );
  OAI222XL U8190 ( .A0(n6379), .A1(n5894), .B0(n2671), .B1(n2661), .C0(n441), 
        .C1(n2662), .Y(n4339) );
  AOI211X1 U8191 ( .A0(n5934), .A1(n2663), .B0(n2672), .C0(n5887), .Y(n2671)
         );
  OAI222XL U8192 ( .A0(n2665), .A1(n5713), .B0(n2666), .B1(n5685), .C0(n6456), 
        .C1(n6506), .Y(n2672) );
  OAI222XL U8193 ( .A0(n6380), .A1(n5894), .B0(n2632), .B1(n2622), .C0(n433), 
        .C1(n2623), .Y(n4331) );
  AOI211X1 U8194 ( .A0(n5934), .A1(n2624), .B0(n2633), .C0(n5887), .Y(n2632)
         );
  OAI222XL U8195 ( .A0(n2626), .A1(n5713), .B0(n2627), .B1(n5685), .C0(n6457), 
        .C1(n5738), .Y(n2633) );
  OAI222XL U8196 ( .A0(n6381), .A1(n5894), .B0(n2593), .B1(n2583), .C0(n425), 
        .C1(n2584), .Y(n4323) );
  AOI211X1 U8197 ( .A0(n5934), .A1(n2585), .B0(n2594), .C0(n5887), .Y(n2593)
         );
  OAI222XL U8198 ( .A0(n2587), .A1(n5713), .B0(n2588), .B1(n5685), .C0(n6458), 
        .C1(n5738), .Y(n2594) );
  OAI222XL U8199 ( .A0(n6382), .A1(n5895), .B0(n2554), .B1(n2544), .C0(n417), 
        .C1(n2545), .Y(n4315) );
  AOI211X1 U8200 ( .A0(n5934), .A1(n2546), .B0(n2555), .C0(n5887), .Y(n2554)
         );
  OAI222XL U8201 ( .A0(n2548), .A1(n5714), .B0(n2549), .B1(n5685), .C0(n6459), 
        .C1(n5738), .Y(n2555) );
  OAI222XL U8202 ( .A0(n6383), .A1(n5895), .B0(n2515), .B1(n2505), .C0(n409), 
        .C1(n2506), .Y(n4307) );
  AOI211X1 U8203 ( .A0(n5934), .A1(n2507), .B0(n2516), .C0(n5887), .Y(n2515)
         );
  OAI222XL U8204 ( .A0(n2509), .A1(n5714), .B0(n2510), .B1(n5685), .C0(n6460), 
        .C1(n5738), .Y(n2516) );
  OAI222XL U8205 ( .A0(n6384), .A1(n5895), .B0(n2476), .B1(n2466), .C0(n401), 
        .C1(n2467), .Y(n4299) );
  AOI211X1 U8206 ( .A0(n5934), .A1(n2468), .B0(n2477), .C0(n5887), .Y(n2476)
         );
  OAI222XL U8207 ( .A0(n2470), .A1(n5714), .B0(n2471), .B1(n5685), .C0(n6461), 
        .C1(n5738), .Y(n2477) );
  OAI222XL U8208 ( .A0(n6385), .A1(n5895), .B0(n2432), .B1(n2422), .C0(n393), 
        .C1(n2423), .Y(n4291) );
  AOI211X1 U8209 ( .A0(n5934), .A1(n2424), .B0(n2433), .C0(n5888), .Y(n2432)
         );
  OAI222XL U8210 ( .A0(n2426), .A1(n5714), .B0(n2427), .B1(n5685), .C0(n6462), 
        .C1(n5738), .Y(n2433) );
  OAI222XL U8211 ( .A0(n6386), .A1(n5895), .B0(n2393), .B1(n2383), .C0(n385), 
        .C1(n2384), .Y(n4283) );
  AOI211X1 U8212 ( .A0(n5934), .A1(n2385), .B0(n2394), .C0(n5888), .Y(n2393)
         );
  OAI222XL U8213 ( .A0(n2387), .A1(n5714), .B0(n2388), .B1(n5685), .C0(n6463), 
        .C1(n5738), .Y(n2394) );
  OAI222XL U8214 ( .A0(n6387), .A1(n5895), .B0(n2354), .B1(n2344), .C0(n377), 
        .C1(n2345), .Y(n4275) );
  AOI211X1 U8215 ( .A0(n5934), .A1(n2346), .B0(n2355), .C0(n5888), .Y(n2354)
         );
  OAI222XL U8216 ( .A0(n2348), .A1(n5714), .B0(n2349), .B1(n5685), .C0(n6464), 
        .C1(n5738), .Y(n2355) );
  OAI222XL U8217 ( .A0(n6388), .A1(n5895), .B0(n2315), .B1(n2305), .C0(n369), 
        .C1(n2306), .Y(n4267) );
  AOI211X1 U8218 ( .A0(n5934), .A1(n2307), .B0(n2316), .C0(n5888), .Y(n2315)
         );
  OAI222XL U8219 ( .A0(n2309), .A1(n5714), .B0(n2310), .B1(n5685), .C0(n6465), 
        .C1(n5738), .Y(n2316) );
  OAI222XL U8220 ( .A0(n6389), .A1(n5895), .B0(n2276), .B1(n2266), .C0(n361), 
        .C1(n2267), .Y(n4259) );
  AOI211X1 U8221 ( .A0(n5934), .A1(n2268), .B0(n2277), .C0(n5888), .Y(n2276)
         );
  OAI222XL U8222 ( .A0(n2270), .A1(n5714), .B0(n2271), .B1(n5685), .C0(n6466), 
        .C1(n5738), .Y(n2277) );
  OAI222XL U8223 ( .A0(n6390), .A1(n5895), .B0(n2237), .B1(n2227), .C0(n353), 
        .C1(n2228), .Y(n4251) );
  AOI211X1 U8224 ( .A0(n5934), .A1(n2229), .B0(n2238), .C0(n5888), .Y(n2237)
         );
  OAI222XL U8225 ( .A0(n2231), .A1(n5714), .B0(n2232), .B1(n5685), .C0(n6467), 
        .C1(n5738), .Y(n2238) );
  OAI222XL U8226 ( .A0(n6391), .A1(n5895), .B0(n2198), .B1(n2188), .C0(n345), 
        .C1(n2189), .Y(n4243) );
  AOI211X1 U8227 ( .A0(n5934), .A1(n2190), .B0(n2199), .C0(n5888), .Y(n2198)
         );
  OAI222XL U8228 ( .A0(n2192), .A1(n5714), .B0(n2193), .B1(n5685), .C0(n6468), 
        .C1(n5738), .Y(n2199) );
  OAI222XL U8229 ( .A0(n6392), .A1(n5895), .B0(n2159), .B1(n2149), .C0(n337), 
        .C1(n2150), .Y(n4235) );
  AOI211X1 U8230 ( .A0(n5934), .A1(n2151), .B0(n2160), .C0(n5888), .Y(n2159)
         );
  OAI222XL U8231 ( .A0(n2153), .A1(n5714), .B0(n2154), .B1(n5685), .C0(n6469), 
        .C1(n5738), .Y(n2160) );
  OAI222XL U8232 ( .A0(n6393), .A1(n5895), .B0(n2115), .B1(n2105), .C0(n329), 
        .C1(n2106), .Y(n4227) );
  AOI211X1 U8233 ( .A0(n5934), .A1(n2107), .B0(n2116), .C0(n5888), .Y(n2115)
         );
  OAI222XL U8234 ( .A0(n2109), .A1(n5714), .B0(n2110), .B1(n5685), .C0(n6470), 
        .C1(n5738), .Y(n2116) );
  OAI222XL U8235 ( .A0(n6394), .A1(n5893), .B0(n2076), .B1(n2066), .C0(n321), 
        .C1(n2067), .Y(n4219) );
  AOI211X1 U8236 ( .A0(n5934), .A1(n2068), .B0(n2077), .C0(n5888), .Y(n2076)
         );
  OAI222XL U8237 ( .A0(n2070), .A1(n5714), .B0(n2071), .B1(n5685), .C0(n6471), 
        .C1(n5738), .Y(n2077) );
  OAI222XL U8238 ( .A0(n6395), .A1(n5894), .B0(n2037), .B1(n2027), .C0(n313), 
        .C1(n2028), .Y(n4211) );
  AOI211X1 U8239 ( .A0(n5934), .A1(n2029), .B0(n2038), .C0(n5888), .Y(n2037)
         );
  OAI222XL U8240 ( .A0(n2031), .A1(n5713), .B0(n2032), .B1(n5684), .C0(n6472), 
        .C1(n5738), .Y(n2038) );
  OAI222XL U8241 ( .A0(n6396), .A1(n5893), .B0(n1996), .B1(n1987), .C0(n305), 
        .C1(n1988), .Y(n4203) );
  AOI211X1 U8242 ( .A0(n5934), .A1(n6473), .B0(n1997), .C0(n5888), .Y(n1996)
         );
  OAI222XL U8243 ( .A0(n1990), .A1(n5714), .B0(n1991), .B1(n5684), .C0(n6474), 
        .C1(n5737), .Y(n1997) );
  OAI222XL U8244 ( .A0(n6397), .A1(n5894), .B0(n1957), .B1(n1948), .C0(n297), 
        .C1(n1949), .Y(n4195) );
  AOI211X1 U8245 ( .A0(n5934), .A1(n6475), .B0(n1958), .C0(n5888), .Y(n1957)
         );
  OAI222XL U8246 ( .A0(n1951), .A1(n5712), .B0(n1952), .B1(n5684), .C0(n6476), 
        .C1(n5737), .Y(n1958) );
  OAI222XL U8247 ( .A0(n6398), .A1(n5895), .B0(n1918), .B1(n1909), .C0(n289), 
        .C1(n1910), .Y(n4187) );
  AOI211X1 U8248 ( .A0(n5934), .A1(n6477), .B0(n1919), .C0(n5889), .Y(n1918)
         );
  OAI222XL U8249 ( .A0(n1912), .A1(n5711), .B0(n1913), .B1(n5684), .C0(n6478), 
        .C1(n5737), .Y(n1919) );
  OAI222XL U8250 ( .A0(n4832), .A1(n5894), .B0(n1879), .B1(n1870), .C0(n281), 
        .C1(n1871), .Y(n4179) );
  AOI211X1 U8251 ( .A0(n5934), .A1(n6479), .B0(n1880), .C0(n5889), .Y(n1879)
         );
  OAI222XL U8252 ( .A0(n1873), .A1(n5711), .B0(n1874), .B1(n5684), .C0(n6480), 
        .C1(n5737), .Y(n1880) );
  OAI222XL U8253 ( .A0(n6399), .A1(n5893), .B0(n1840), .B1(n1831), .C0(n273), 
        .C1(n4643), .Y(n4171) );
  AOI211X1 U8254 ( .A0(n5934), .A1(n6481), .B0(n1841), .C0(n5889), .Y(n1840)
         );
  OAI222XL U8255 ( .A0(n1834), .A1(n5711), .B0(n1835), .B1(n5684), .C0(n6482), 
        .C1(n5737), .Y(n1841) );
  OAI222XL U8256 ( .A0(n1790), .A1(n5712), .B0(n1791), .B1(n5684), .C0(n6484), 
        .C1(n5737), .Y(n1797) );
  OAI222XL U8257 ( .A0(n1745), .A1(n5714), .B0(n1746), .B1(n5684), .C0(n6486), 
        .C1(n5737), .Y(n1752) );
  OAI222XL U8258 ( .A0(n6402), .A1(n5893), .B0(n1707), .B1(n1698), .C0(n249), 
        .C1(n1699), .Y(n4147) );
  AOI211X1 U8259 ( .A0(n5934), .A1(n6487), .B0(n1708), .C0(n5889), .Y(n1707)
         );
  OAI222XL U8260 ( .A0(n1701), .A1(n5711), .B0(n1702), .B1(n5684), .C0(n6488), 
        .C1(n5737), .Y(n1708) );
  OAI222XL U8261 ( .A0(n6403), .A1(n5895), .B0(n1663), .B1(n1654), .C0(n241), 
        .C1(n1655), .Y(n4139) );
  AOI211X1 U8262 ( .A0(n5934), .A1(n6489), .B0(n1664), .C0(n5889), .Y(n1663)
         );
  OAI222XL U8263 ( .A0(n1657), .A1(n5713), .B0(n1658), .B1(n5684), .C0(n6490), 
        .C1(n5737), .Y(n1664) );
  OAI222XL U8264 ( .A0(n6404), .A1(n5895), .B0(n1619), .B1(n1610), .C0(n233), 
        .C1(n1611), .Y(n4131) );
  AOI211X1 U8265 ( .A0(n5934), .A1(n6491), .B0(n1620), .C0(n5889), .Y(n1619)
         );
  OAI222XL U8266 ( .A0(n1613), .A1(n5712), .B0(n1614), .B1(n5684), .C0(n6492), 
        .C1(n5737), .Y(n1620) );
  OAI222XL U8267 ( .A0(n6405), .A1(n5894), .B0(n1575), .B1(n1566), .C0(n225), 
        .C1(n1567), .Y(n4123) );
  AOI211X1 U8268 ( .A0(n5934), .A1(n6493), .B0(n1576), .C0(n5889), .Y(n1575)
         );
  OAI222XL U8269 ( .A0(n1569), .A1(n5714), .B0(n1570), .B1(n5684), .C0(n6494), 
        .C1(n5737), .Y(n1576) );
  OAI222XL U8270 ( .A0(n6406), .A1(n5895), .B0(n1531), .B1(n1522), .C0(n217), 
        .C1(n1523), .Y(n4115) );
  AOI211X1 U8271 ( .A0(n5934), .A1(n6495), .B0(n1532), .C0(n5889), .Y(n1531)
         );
  OAI222XL U8272 ( .A0(n1525), .A1(n5712), .B0(n1526), .B1(n5684), .C0(n6496), 
        .C1(n5737), .Y(n1532) );
  OAI222XL U8273 ( .A0(n6407), .A1(n5893), .B0(n1487), .B1(n1478), .C0(n209), 
        .C1(n1479), .Y(n4107) );
  AOI211X1 U8274 ( .A0(n5935), .A1(n6497), .B0(n1488), .C0(n5889), .Y(n1487)
         );
  OAI222XL U8275 ( .A0(n1481), .A1(n5713), .B0(n1482), .B1(n5686), .C0(n6498), 
        .C1(n5738), .Y(n1488) );
  OAI222XL U8276 ( .A0(n6347), .A1(n5903), .B0(n3937), .B1(n3929), .C0(n696), 
        .C1(n3930), .Y(n4594) );
  AOI211X1 U8277 ( .A0(n5941), .A1(n3931), .B0(n3938), .C0(n5896), .Y(n3937)
         );
  OAI222XL U8278 ( .A0(n3933), .A1(n5708), .B0(n3934), .B1(n5682), .C0(n6424), 
        .C1(n6505), .Y(n3938) );
  OAI222XL U8279 ( .A0(n6348), .A1(n5903), .B0(n3898), .B1(n3890), .C0(n688), 
        .C1(n3891), .Y(n4586) );
  AOI211X1 U8280 ( .A0(n5941), .A1(n3892), .B0(n3899), .C0(n5896), .Y(n3898)
         );
  OAI222XL U8281 ( .A0(n3894), .A1(n5708), .B0(n3895), .B1(n5683), .C0(n6425), 
        .C1(n5736), .Y(n3899) );
  OAI222XL U8282 ( .A0(n6349), .A1(n5903), .B0(n3859), .B1(n3851), .C0(n680), 
        .C1(n3852), .Y(n4578) );
  AOI211X1 U8283 ( .A0(n5941), .A1(n3853), .B0(n3860), .C0(n5896), .Y(n3859)
         );
  OAI222XL U8284 ( .A0(n3855), .A1(n5710), .B0(n3856), .B1(n5683), .C0(n6426), 
        .C1(n5734), .Y(n3860) );
  OAI222XL U8285 ( .A0(n6350), .A1(n5903), .B0(n3820), .B1(n3812), .C0(n672), 
        .C1(n3813), .Y(n4570) );
  AOI211X1 U8286 ( .A0(n5941), .A1(n3814), .B0(n3821), .C0(n5896), .Y(n3820)
         );
  OAI222XL U8287 ( .A0(n3816), .A1(n5710), .B0(n3817), .B1(n5683), .C0(n6427), 
        .C1(n5734), .Y(n3821) );
  OAI222XL U8288 ( .A0(n6351), .A1(n5903), .B0(n3781), .B1(n3773), .C0(n664), 
        .C1(n3774), .Y(n4562) );
  AOI211X1 U8289 ( .A0(n5941), .A1(n3775), .B0(n3782), .C0(n5896), .Y(n3781)
         );
  OAI222XL U8290 ( .A0(n3777), .A1(n5709), .B0(n3778), .B1(n5683), .C0(n6428), 
        .C1(n6505), .Y(n3782) );
  OAI222XL U8291 ( .A0(n6352), .A1(n5903), .B0(n3742), .B1(n3734), .C0(n656), 
        .C1(n3735), .Y(n4554) );
  AOI211X1 U8292 ( .A0(n5941), .A1(n3736), .B0(n3743), .C0(n5896), .Y(n3742)
         );
  OAI222XL U8293 ( .A0(n3738), .A1(n5708), .B0(n3739), .B1(n5683), .C0(n6429), 
        .C1(n5736), .Y(n3743) );
  OAI222XL U8294 ( .A0(n6353), .A1(n5903), .B0(n3698), .B1(n3690), .C0(n648), 
        .C1(n5670), .Y(n4546) );
  AOI211X1 U8295 ( .A0(n5941), .A1(n3692), .B0(n3699), .C0(n5896), .Y(n3698)
         );
  OAI222XL U8296 ( .A0(n3694), .A1(n6500), .B0(n3695), .B1(n5683), .C0(n6430), 
        .C1(n6505), .Y(n3699) );
  OAI222XL U8297 ( .A0(n6354), .A1(n5903), .B0(n3659), .B1(n3651), .C0(n640), 
        .C1(n3652), .Y(n4538) );
  AOI211X1 U8298 ( .A0(n5941), .A1(n3653), .B0(n3660), .C0(n5896), .Y(n3659)
         );
  OAI222XL U8299 ( .A0(n3655), .A1(n5709), .B0(n3656), .B1(n5683), .C0(n6431), 
        .C1(n6505), .Y(n3660) );
  OAI222XL U8300 ( .A0(n6355), .A1(n5903), .B0(n3620), .B1(n3612), .C0(n632), 
        .C1(n3613), .Y(n4530) );
  AOI211X1 U8301 ( .A0(n5941), .A1(n3614), .B0(n3621), .C0(n5896), .Y(n3620)
         );
  OAI222XL U8302 ( .A0(n3616), .A1(n5710), .B0(n3617), .B1(n5683), .C0(n6432), 
        .C1(n5733), .Y(n3621) );
  OAI222XL U8303 ( .A0(n6356), .A1(n5903), .B0(n3581), .B1(n3573), .C0(n624), 
        .C1(n3574), .Y(n4522) );
  AOI211X1 U8304 ( .A0(n5941), .A1(n3575), .B0(n3582), .C0(n5896), .Y(n3581)
         );
  OAI222XL U8305 ( .A0(n3577), .A1(n5709), .B0(n3578), .B1(n5683), .C0(n6433), 
        .C1(n5736), .Y(n3582) );
  OAI222XL U8306 ( .A0(n6357), .A1(n5903), .B0(n3542), .B1(n3534), .C0(n616), 
        .C1(n3535), .Y(n4514) );
  AOI211X1 U8307 ( .A0(n5941), .A1(n3536), .B0(n3543), .C0(n5896), .Y(n3542)
         );
  OAI222XL U8308 ( .A0(n3538), .A1(n6500), .B0(n3539), .B1(n5683), .C0(n6434), 
        .C1(n5735), .Y(n3543) );
  OAI222XL U8309 ( .A0(n6358), .A1(n5905), .B0(n3503), .B1(n3495), .C0(n608), 
        .C1(n3496), .Y(n4506) );
  AOI211X1 U8310 ( .A0(n5941), .A1(n3497), .B0(n3504), .C0(n5896), .Y(n3503)
         );
  OAI222XL U8311 ( .A0(n3499), .A1(n5708), .B0(n3500), .B1(n5683), .C0(n6435), 
        .C1(n5734), .Y(n3504) );
  OAI222XL U8312 ( .A0(n6359), .A1(n5904), .B0(n3464), .B1(n3456), .C0(n600), 
        .C1(n3457), .Y(n4498) );
  AOI211X1 U8313 ( .A0(n5941), .A1(n3458), .B0(n3465), .C0(n5897), .Y(n3464)
         );
  OAI222XL U8314 ( .A0(n3460), .A1(n5708), .B0(n3461), .B1(n5683), .C0(n6436), 
        .C1(n5734), .Y(n3465) );
  OAI222XL U8315 ( .A0(n6360), .A1(n5903), .B0(n3425), .B1(n3417), .C0(n592), 
        .C1(n3418), .Y(n4490) );
  AOI211X1 U8316 ( .A0(n5941), .A1(n3419), .B0(n3426), .C0(n5897), .Y(n3425)
         );
  OAI222XL U8317 ( .A0(n3421), .A1(n5708), .B0(n3422), .B1(n5683), .C0(n6437), 
        .C1(n5734), .Y(n3426) );
  OAI222XL U8318 ( .A0(n6361), .A1(n5905), .B0(n3381), .B1(n3373), .C0(n584), 
        .C1(n3374), .Y(n4482) );
  AOI211X1 U8319 ( .A0(n5941), .A1(n3375), .B0(n3382), .C0(n5897), .Y(n3381)
         );
  OAI222XL U8320 ( .A0(n3377), .A1(n5708), .B0(n3378), .B1(n5683), .C0(n6438), 
        .C1(n6505), .Y(n3382) );
  OAI222XL U8321 ( .A0(n6362), .A1(n5904), .B0(n3342), .B1(n3334), .C0(n576), 
        .C1(n3335), .Y(n4474) );
  AOI211X1 U8322 ( .A0(n5941), .A1(n3336), .B0(n3343), .C0(n5897), .Y(n3342)
         );
  OAI222XL U8323 ( .A0(n3338), .A1(n5708), .B0(n3339), .B1(n5683), .C0(n6439), 
        .C1(n5734), .Y(n3343) );
  OAI222XL U8324 ( .A0(n6363), .A1(n5903), .B0(n3303), .B1(n3295), .C0(n568), 
        .C1(n3296), .Y(n4466) );
  AOI211X1 U8325 ( .A0(n5941), .A1(n3297), .B0(n3304), .C0(n5897), .Y(n3303)
         );
  OAI222XL U8326 ( .A0(n3299), .A1(n5708), .B0(n3300), .B1(n5683), .C0(n6440), 
        .C1(n6505), .Y(n3304) );
  OAI222XL U8327 ( .A0(n6364), .A1(n5905), .B0(n3264), .B1(n3256), .C0(n560), 
        .C1(n3257), .Y(n4458) );
  AOI211X1 U8328 ( .A0(n5941), .A1(n3258), .B0(n3265), .C0(n5897), .Y(n3264)
         );
  OAI222XL U8329 ( .A0(n3260), .A1(n5708), .B0(n3261), .B1(n6418), .C0(n6441), 
        .C1(n5734), .Y(n3265) );
  OAI222XL U8330 ( .A0(n6365), .A1(n5904), .B0(n3225), .B1(n3217), .C0(n552), 
        .C1(n3218), .Y(n4450) );
  AOI211X1 U8331 ( .A0(n5941), .A1(n3219), .B0(n3226), .C0(n5897), .Y(n3225)
         );
  OAI222XL U8332 ( .A0(n3221), .A1(n5708), .B0(n3222), .B1(n5682), .C0(n6442), 
        .C1(n5736), .Y(n3226) );
  OAI222XL U8333 ( .A0(n6366), .A1(n5903), .B0(n3186), .B1(n3178), .C0(n544), 
        .C1(n3179), .Y(n4442) );
  AOI211X1 U8334 ( .A0(n5941), .A1(n3180), .B0(n3187), .C0(n5897), .Y(n3186)
         );
  OAI222XL U8335 ( .A0(n3182), .A1(n5708), .B0(n3183), .B1(n5683), .C0(n6443), 
        .C1(n5736), .Y(n3187) );
  OAI222XL U8336 ( .A0(n6367), .A1(n5903), .B0(n3147), .B1(n3139), .C0(n536), 
        .C1(n4674), .Y(n4434) );
  AOI211X1 U8337 ( .A0(n5941), .A1(n3141), .B0(n3148), .C0(n5897), .Y(n3147)
         );
  OAI222XL U8338 ( .A0(n3143), .A1(n5708), .B0(n3144), .B1(n5683), .C0(n6444), 
        .C1(n5736), .Y(n3148) );
  OAI222XL U8339 ( .A0(n6368), .A1(n5905), .B0(n3108), .B1(n3100), .C0(n528), 
        .C1(n3101), .Y(n4426) );
  AOI211X1 U8340 ( .A0(n5941), .A1(n3102), .B0(n3109), .C0(n5897), .Y(n3108)
         );
  OAI222XL U8341 ( .A0(n3104), .A1(n5708), .B0(n3105), .B1(n5681), .C0(n6445), 
        .C1(n5736), .Y(n3109) );
  OAI222XL U8342 ( .A0(n6369), .A1(n5904), .B0(n3064), .B1(n3056), .C0(n520), 
        .C1(n3057), .Y(n4418) );
  AOI211X1 U8343 ( .A0(n5941), .A1(n3058), .B0(n3065), .C0(n5897), .Y(n3064)
         );
  OAI222XL U8344 ( .A0(n3060), .A1(n5708), .B0(n3061), .B1(n5683), .C0(n6446), 
        .C1(n5736), .Y(n3065) );
  OAI222XL U8345 ( .A0(n6370), .A1(n5904), .B0(n3025), .B1(n3017), .C0(n512), 
        .C1(n3018), .Y(n4410) );
  AOI211X1 U8346 ( .A0(n5941), .A1(n3019), .B0(n3026), .C0(n5897), .Y(n3025)
         );
  OAI222XL U8347 ( .A0(n3021), .A1(n5709), .B0(n3022), .B1(n5681), .C0(n6447), 
        .C1(n5736), .Y(n3026) );
  OAI222XL U8348 ( .A0(n6371), .A1(n5904), .B0(n2986), .B1(n2978), .C0(n504), 
        .C1(n2979), .Y(n4402) );
  AOI211X1 U8349 ( .A0(n5941), .A1(n2980), .B0(n2987), .C0(n5897), .Y(n2986)
         );
  OAI222XL U8350 ( .A0(n2982), .A1(n5709), .B0(n2983), .B1(n5683), .C0(n6448), 
        .C1(n5736), .Y(n2987) );
  OAI222XL U8351 ( .A0(n6372), .A1(n5904), .B0(n2947), .B1(n2939), .C0(n496), 
        .C1(n4675), .Y(n4394) );
  AOI211X1 U8352 ( .A0(n5941), .A1(n2941), .B0(n2948), .C0(n5898), .Y(n2947)
         );
  OAI222XL U8353 ( .A0(n2943), .A1(n5709), .B0(n2944), .B1(n5682), .C0(n6449), 
        .C1(n5736), .Y(n2948) );
  OAI222XL U8354 ( .A0(n6373), .A1(n5904), .B0(n2908), .B1(n2900), .C0(n488), 
        .C1(n2901), .Y(n4386) );
  AOI211X1 U8355 ( .A0(n5941), .A1(n2902), .B0(n2909), .C0(n5898), .Y(n2908)
         );
  OAI222XL U8356 ( .A0(n2904), .A1(n5709), .B0(n2905), .B1(n6418), .C0(n6450), 
        .C1(n5736), .Y(n2909) );
  OAI222XL U8357 ( .A0(n6374), .A1(n5904), .B0(n2869), .B1(n2861), .C0(n480), 
        .C1(n2862), .Y(n4378) );
  AOI211X1 U8358 ( .A0(n5941), .A1(n2863), .B0(n2870), .C0(n5898), .Y(n2869)
         );
  OAI222XL U8359 ( .A0(n2865), .A1(n5709), .B0(n2866), .B1(n5683), .C0(n6451), 
        .C1(n5736), .Y(n2870) );
  OAI222XL U8360 ( .A0(n6375), .A1(n5904), .B0(n2830), .B1(n2822), .C0(n472), 
        .C1(n2823), .Y(n4370) );
  AOI211X1 U8361 ( .A0(n5941), .A1(n2824), .B0(n2831), .C0(n5898), .Y(n2830)
         );
  OAI222XL U8362 ( .A0(n2826), .A1(n5709), .B0(n2827), .B1(n6418), .C0(n6452), 
        .C1(n5736), .Y(n2831) );
  OAI222XL U8363 ( .A0(n6376), .A1(n5904), .B0(n2791), .B1(n2783), .C0(n464), 
        .C1(n2784), .Y(n4362) );
  AOI211X1 U8364 ( .A0(n5940), .A1(n2785), .B0(n2792), .C0(n5898), .Y(n2791)
         );
  OAI222XL U8365 ( .A0(n2787), .A1(n5709), .B0(n2788), .B1(n6418), .C0(n6453), 
        .C1(n5736), .Y(n2792) );
  OAI222XL U8366 ( .A0(n6377), .A1(n5904), .B0(n2747), .B1(n2739), .C0(n456), 
        .C1(n2740), .Y(n4354) );
  AOI211X1 U8367 ( .A0(n5940), .A1(n2741), .B0(n2748), .C0(n5898), .Y(n2747)
         );
  OAI222XL U8368 ( .A0(n2743), .A1(n5709), .B0(n2744), .B1(n6418), .C0(n6454), 
        .C1(n5736), .Y(n2748) );
  OAI222XL U8369 ( .A0(n6378), .A1(n5904), .B0(n2708), .B1(n2700), .C0(n448), 
        .C1(n2701), .Y(n4346) );
  AOI211X1 U8370 ( .A0(n5940), .A1(n2702), .B0(n2709), .C0(n5898), .Y(n2708)
         );
  OAI222XL U8371 ( .A0(n2704), .A1(n5709), .B0(n2705), .B1(n6418), .C0(n6455), 
        .C1(n5736), .Y(n2709) );
  OAI222XL U8372 ( .A0(n6379), .A1(n5904), .B0(n2669), .B1(n2661), .C0(n440), 
        .C1(n2662), .Y(n4338) );
  AOI211X1 U8373 ( .A0(n5940), .A1(n2663), .B0(n2670), .C0(n5898), .Y(n2669)
         );
  OAI222XL U8374 ( .A0(n2665), .A1(n5709), .B0(n2666), .B1(n5682), .C0(n6456), 
        .C1(n5736), .Y(n2670) );
  OAI222XL U8375 ( .A0(n6380), .A1(n5904), .B0(n2630), .B1(n2622), .C0(n432), 
        .C1(n2623), .Y(n4330) );
  AOI211X1 U8376 ( .A0(n5940), .A1(n2624), .B0(n2631), .C0(n5898), .Y(n2630)
         );
  OAI222XL U8377 ( .A0(n2626), .A1(n5709), .B0(n2627), .B1(n5682), .C0(n6457), 
        .C1(n5733), .Y(n2631) );
  OAI222XL U8378 ( .A0(n6381), .A1(n5904), .B0(n2591), .B1(n2583), .C0(n424), 
        .C1(n2584), .Y(n4322) );
  AOI211X1 U8379 ( .A0(n5940), .A1(n2585), .B0(n2592), .C0(n5898), .Y(n2591)
         );
  OAI222XL U8380 ( .A0(n2587), .A1(n5709), .B0(n2588), .B1(n5682), .C0(n6458), 
        .C1(n5733), .Y(n2592) );
  OAI222XL U8381 ( .A0(n6382), .A1(n5905), .B0(n2552), .B1(n2544), .C0(n416), 
        .C1(n2545), .Y(n4314) );
  AOI211X1 U8382 ( .A0(n5940), .A1(n2546), .B0(n2553), .C0(n5898), .Y(n2552)
         );
  OAI222XL U8383 ( .A0(n2548), .A1(n5710), .B0(n2549), .B1(n5682), .C0(n6459), 
        .C1(n5733), .Y(n2553) );
  OAI222XL U8384 ( .A0(n6383), .A1(n5905), .B0(n2513), .B1(n2505), .C0(n408), 
        .C1(n2506), .Y(n4306) );
  AOI211X1 U8385 ( .A0(n5940), .A1(n2507), .B0(n2514), .C0(n5898), .Y(n2513)
         );
  OAI222XL U8386 ( .A0(n2509), .A1(n5710), .B0(n2510), .B1(n5682), .C0(n6460), 
        .C1(n5733), .Y(n2514) );
  OAI222XL U8387 ( .A0(n6384), .A1(n5905), .B0(n2474), .B1(n2466), .C0(n400), 
        .C1(n2467), .Y(n4298) );
  AOI211X1 U8388 ( .A0(n5940), .A1(n2468), .B0(n2475), .C0(n5898), .Y(n2474)
         );
  OAI222XL U8389 ( .A0(n2470), .A1(n5710), .B0(n2471), .B1(n5682), .C0(n6461), 
        .C1(n5733), .Y(n2475) );
  OAI222XL U8390 ( .A0(n6385), .A1(n5905), .B0(n2430), .B1(n2422), .C0(n392), 
        .C1(n2423), .Y(n4290) );
  AOI211X1 U8391 ( .A0(n5940), .A1(n2424), .B0(n2431), .C0(n4647), .Y(n2430)
         );
  OAI222XL U8392 ( .A0(n2426), .A1(n5710), .B0(n2427), .B1(n5682), .C0(n6462), 
        .C1(n5733), .Y(n2431) );
  OAI222XL U8393 ( .A0(n6386), .A1(n5905), .B0(n2391), .B1(n2383), .C0(n384), 
        .C1(n2384), .Y(n4282) );
  AOI211X1 U8394 ( .A0(n5940), .A1(n2385), .B0(n2392), .C0(n4647), .Y(n2391)
         );
  OAI222XL U8395 ( .A0(n2387), .A1(n5710), .B0(n2388), .B1(n5682), .C0(n6463), 
        .C1(n5733), .Y(n2392) );
  OAI222XL U8396 ( .A0(n6387), .A1(n5905), .B0(n2352), .B1(n2344), .C0(n376), 
        .C1(n2345), .Y(n4274) );
  AOI211X1 U8397 ( .A0(n5940), .A1(n2346), .B0(n2353), .C0(n4647), .Y(n2352)
         );
  OAI222XL U8398 ( .A0(n2348), .A1(n5710), .B0(n2349), .B1(n5682), .C0(n6464), 
        .C1(n5733), .Y(n2353) );
  OAI222XL U8399 ( .A0(n6388), .A1(n5905), .B0(n2313), .B1(n2305), .C0(n368), 
        .C1(n2306), .Y(n4266) );
  AOI211X1 U8400 ( .A0(n5940), .A1(n2307), .B0(n2314), .C0(n5896), .Y(n2313)
         );
  OAI222XL U8401 ( .A0(n2309), .A1(n5710), .B0(n2310), .B1(n5682), .C0(n6465), 
        .C1(n5733), .Y(n2314) );
  OAI222XL U8402 ( .A0(n6389), .A1(n5905), .B0(n2274), .B1(n2266), .C0(n360), 
        .C1(n2267), .Y(n4258) );
  AOI211X1 U8403 ( .A0(n5940), .A1(n2268), .B0(n2275), .C0(n4647), .Y(n2274)
         );
  OAI222XL U8404 ( .A0(n2270), .A1(n5710), .B0(n2271), .B1(n5682), .C0(n6466), 
        .C1(n5733), .Y(n2275) );
  OAI222XL U8405 ( .A0(n6390), .A1(n5905), .B0(n2235), .B1(n2227), .C0(n352), 
        .C1(n2228), .Y(n4250) );
  AOI211X1 U8406 ( .A0(n5940), .A1(n2229), .B0(n2236), .C0(n5896), .Y(n2235)
         );
  OAI222XL U8407 ( .A0(n2231), .A1(n5710), .B0(n2232), .B1(n5682), .C0(n6467), 
        .C1(n5733), .Y(n2236) );
  OAI222XL U8408 ( .A0(n6391), .A1(n5905), .B0(n2196), .B1(n2188), .C0(n344), 
        .C1(n2189), .Y(n4242) );
  AOI211X1 U8409 ( .A0(n5940), .A1(n2190), .B0(n2197), .C0(n4647), .Y(n2196)
         );
  OAI222XL U8410 ( .A0(n2192), .A1(n5710), .B0(n2193), .B1(n5682), .C0(n6468), 
        .C1(n5736), .Y(n2197) );
  OAI222XL U8411 ( .A0(n6392), .A1(n5905), .B0(n2157), .B1(n2149), .C0(n336), 
        .C1(n2150), .Y(n4234) );
  AOI211X1 U8412 ( .A0(n5940), .A1(n2151), .B0(n2158), .C0(n4647), .Y(n2157)
         );
  OAI222XL U8413 ( .A0(n2153), .A1(n5710), .B0(n2154), .B1(n5682), .C0(n6469), 
        .C1(n5734), .Y(n2158) );
  OAI222XL U8414 ( .A0(n6393), .A1(n5905), .B0(n2113), .B1(n2105), .C0(n328), 
        .C1(n2106), .Y(n4226) );
  AOI211X1 U8415 ( .A0(n5940), .A1(n2107), .B0(n2114), .C0(n5896), .Y(n2113)
         );
  OAI222XL U8416 ( .A0(n2109), .A1(n5710), .B0(n2110), .B1(n5682), .C0(n6470), 
        .C1(n5736), .Y(n2114) );
  OAI222XL U8417 ( .A0(n6394), .A1(n5903), .B0(n2074), .B1(n2066), .C0(n320), 
        .C1(n2067), .Y(n4218) );
  AOI211X1 U8418 ( .A0(n5940), .A1(n2068), .B0(n2075), .C0(n4647), .Y(n2074)
         );
  OAI222XL U8419 ( .A0(n2070), .A1(n5708), .B0(n2071), .B1(n5682), .C0(n6471), 
        .C1(n5733), .Y(n2075) );
  OAI222XL U8420 ( .A0(n6395), .A1(n5903), .B0(n2035), .B1(n2027), .C0(n312), 
        .C1(n2028), .Y(n4210) );
  AOI211X1 U8421 ( .A0(n5940), .A1(n2029), .B0(n2036), .C0(n5896), .Y(n2035)
         );
  OAI222XL U8422 ( .A0(n2031), .A1(n5709), .B0(n2032), .B1(n5681), .C0(n6472), 
        .C1(n5734), .Y(n2036) );
  OAI222XL U8423 ( .A0(n6396), .A1(n5905), .B0(n1994), .B1(n1987), .C0(n304), 
        .C1(n1988), .Y(n4202) );
  AOI211X1 U8424 ( .A0(n5940), .A1(n6473), .B0(n1995), .C0(n5896), .Y(n1994)
         );
  OAI222XL U8425 ( .A0(n1990), .A1(n5708), .B0(n1991), .B1(n5681), .C0(n6474), 
        .C1(n5735), .Y(n1995) );
  OAI222XL U8426 ( .A0(n6397), .A1(n5905), .B0(n1955), .B1(n1948), .C0(n296), 
        .C1(n1949), .Y(n4194) );
  AOI211X1 U8427 ( .A0(n5940), .A1(n6475), .B0(n1956), .C0(n4647), .Y(n1955)
         );
  OAI222XL U8428 ( .A0(n1951), .A1(n5710), .B0(n1952), .B1(n5681), .C0(n6476), 
        .C1(n5735), .Y(n1956) );
  OAI222XL U8429 ( .A0(n6398), .A1(n5905), .B0(n1916), .B1(n1909), .C0(n288), 
        .C1(n1910), .Y(n4186) );
  AOI211X1 U8430 ( .A0(n5940), .A1(n6477), .B0(n1917), .C0(n4647), .Y(n1916)
         );
  OAI222XL U8431 ( .A0(n1912), .A1(n5710), .B0(n1913), .B1(n5681), .C0(n6478), 
        .C1(n5735), .Y(n1917) );
  OAI222XL U8432 ( .A0(n4832), .A1(n5904), .B0(n1877), .B1(n1870), .C0(n280), 
        .C1(n1871), .Y(n4178) );
  AOI211X1 U8433 ( .A0(n5940), .A1(n6479), .B0(n1878), .C0(n4647), .Y(n1877)
         );
  OAI222XL U8434 ( .A0(n1873), .A1(n5710), .B0(n1874), .B1(n5681), .C0(n6480), 
        .C1(n5735), .Y(n1878) );
  OAI222XL U8435 ( .A0(n6399), .A1(n5904), .B0(n1838), .B1(n1831), .C0(n272), 
        .C1(n4643), .Y(n4170) );
  AOI211X1 U8436 ( .A0(n5940), .A1(n6481), .B0(n1839), .C0(n4647), .Y(n1838)
         );
  OAI222XL U8437 ( .A0(n1834), .A1(n5709), .B0(n1835), .B1(n5681), .C0(n6482), 
        .C1(n5735), .Y(n1839) );
  OAI222XL U8438 ( .A0(n6400), .A1(n5904), .B0(n1794), .B1(n1787), .C0(n264), 
        .C1(n1788), .Y(n4162) );
  AOI211X1 U8439 ( .A0(n5940), .A1(n6483), .B0(n1795), .C0(n4647), .Y(n1794)
         );
  OAI222XL U8440 ( .A0(n1790), .A1(n5708), .B0(n1791), .B1(n5681), .C0(n6484), 
        .C1(n5735), .Y(n1795) );
  OAI222XL U8441 ( .A0(n6401), .A1(n5903), .B0(n1749), .B1(n1742), .C0(n256), 
        .C1(n1743), .Y(n4154) );
  AOI211X1 U8442 ( .A0(n5940), .A1(n6485), .B0(n1750), .C0(n4647), .Y(n1749)
         );
  OAI222XL U8443 ( .A0(n1745), .A1(n5709), .B0(n1746), .B1(n5681), .C0(n6486), 
        .C1(n5735), .Y(n1750) );
  OAI222XL U8444 ( .A0(n6402), .A1(n5905), .B0(n1705), .B1(n1698), .C0(n248), 
        .C1(n1699), .Y(n4146) );
  AOI211X1 U8445 ( .A0(n5940), .A1(n6487), .B0(n1706), .C0(n4647), .Y(n1705)
         );
  OAI222XL U8446 ( .A0(n1701), .A1(n5708), .B0(n1702), .B1(n5681), .C0(n6488), 
        .C1(n5735), .Y(n1706) );
  OAI222XL U8447 ( .A0(n6403), .A1(n5904), .B0(n1661), .B1(n1654), .C0(n240), 
        .C1(n1655), .Y(n4138) );
  AOI211X1 U8448 ( .A0(n5940), .A1(n6489), .B0(n1662), .C0(n4647), .Y(n1661)
         );
  OAI222XL U8449 ( .A0(n1657), .A1(n5709), .B0(n1658), .B1(n5681), .C0(n6490), 
        .C1(n5735), .Y(n1662) );
  OAI222XL U8450 ( .A0(n6404), .A1(n5904), .B0(n1617), .B1(n1610), .C0(n232), 
        .C1(n1611), .Y(n4130) );
  AOI211X1 U8451 ( .A0(n5940), .A1(n6491), .B0(n1618), .C0(n4647), .Y(n1617)
         );
  OAI222XL U8452 ( .A0(n1613), .A1(n5710), .B0(n1614), .B1(n5681), .C0(n6492), 
        .C1(n5735), .Y(n1618) );
  OAI222XL U8453 ( .A0(n6405), .A1(n5903), .B0(n1573), .B1(n1566), .C0(n224), 
        .C1(n1567), .Y(n4122) );
  AOI211X1 U8454 ( .A0(n5940), .A1(n6493), .B0(n1574), .C0(n4647), .Y(n1573)
         );
  OAI222XL U8455 ( .A0(n1569), .A1(n5709), .B0(n1570), .B1(n5681), .C0(n6494), 
        .C1(n5735), .Y(n1574) );
  OAI222XL U8456 ( .A0(n6406), .A1(n5903), .B0(n1529), .B1(n1522), .C0(n216), 
        .C1(n1523), .Y(n4114) );
  AOI211X1 U8457 ( .A0(n5940), .A1(n6495), .B0(n1530), .C0(n4647), .Y(n1529)
         );
  OAI222XL U8458 ( .A0(n1525), .A1(n6500), .B0(n1526), .B1(n5681), .C0(n6496), 
        .C1(n5735), .Y(n1530) );
  OAI222XL U8459 ( .A0(n6407), .A1(n5905), .B0(n1485), .B1(n1478), .C0(n208), 
        .C1(n1479), .Y(n4106) );
  AOI211X1 U8460 ( .A0(n5941), .A1(n6497), .B0(n1486), .C0(n4647), .Y(n1485)
         );
  OAI222XL U8461 ( .A0(n1481), .A1(n5710), .B0(n1482), .B1(n5682), .C0(n6498), 
        .C1(n5736), .Y(n1486) );
  OAI222XL U8462 ( .A0(n6347), .A1(n5909), .B0(n3928), .B1(n3929), .C0(n694), 
        .C1(n3930), .Y(n4592) );
  AOI211X1 U8463 ( .A0(n5948), .A1(n3931), .B0(n3932), .C0(n5760), .Y(n3928)
         );
  OAI222XL U8464 ( .A0(n3933), .A1(n5702), .B0(n3934), .B1(n5676), .C0(n6424), 
        .C1(n6260), .Y(n3932) );
  OAI222XL U8465 ( .A0(n6348), .A1(n5909), .B0(n3889), .B1(n3890), .C0(n686), 
        .C1(n3891), .Y(n4584) );
  AOI211X1 U8466 ( .A0(n5948), .A1(n3892), .B0(n3893), .C0(n5758), .Y(n3889)
         );
  OAI222XL U8467 ( .A0(n3894), .A1(n5702), .B0(n3895), .B1(n5677), .C0(n6425), 
        .C1(n5729), .Y(n3893) );
  OAI222XL U8468 ( .A0(n6349), .A1(n5909), .B0(n3850), .B1(n3851), .C0(n678), 
        .C1(n3852), .Y(n4576) );
  AOI211X1 U8469 ( .A0(n5948), .A1(n3853), .B0(n3854), .C0(n5759), .Y(n3850)
         );
  OAI222XL U8470 ( .A0(n3855), .A1(n5702), .B0(n3856), .B1(n5677), .C0(n6426), 
        .C1(n6503), .Y(n3854) );
  OAI222XL U8471 ( .A0(n6350), .A1(n5909), .B0(n3811), .B1(n3812), .C0(n670), 
        .C1(n3813), .Y(n4568) );
  AOI211X1 U8472 ( .A0(n5948), .A1(n3814), .B0(n3815), .C0(n5758), .Y(n3811)
         );
  OAI222XL U8473 ( .A0(n3816), .A1(n5703), .B0(n3817), .B1(n5677), .C0(n6427), 
        .C1(n6503), .Y(n3815) );
  OAI222XL U8474 ( .A0(n6351), .A1(n5909), .B0(n3772), .B1(n3773), .C0(n662), 
        .C1(n3774), .Y(n4560) );
  AOI211X1 U8475 ( .A0(n5948), .A1(n3775), .B0(n3776), .C0(n5760), .Y(n3772)
         );
  OAI222XL U8476 ( .A0(n3777), .A1(n5702), .B0(n3778), .B1(n5677), .C0(n6428), 
        .C1(n6503), .Y(n3776) );
  OAI222XL U8477 ( .A0(n6352), .A1(n5909), .B0(n3733), .B1(n3734), .C0(n654), 
        .C1(n3735), .Y(n4552) );
  AOI211X1 U8478 ( .A0(n5948), .A1(n3736), .B0(n3737), .C0(n5758), .Y(n3733)
         );
  OAI222XL U8479 ( .A0(n3738), .A1(n5703), .B0(n3739), .B1(n5677), .C0(n6429), 
        .C1(n5729), .Y(n3737) );
  OAI222XL U8480 ( .A0(n6353), .A1(n5909), .B0(n3689), .B1(n3690), .C0(n646), 
        .C1(n5670), .Y(n4544) );
  AOI211X1 U8481 ( .A0(n5948), .A1(n3692), .B0(n3693), .C0(n5759), .Y(n3689)
         );
  OAI222XL U8482 ( .A0(n3694), .A1(n5704), .B0(n3695), .B1(n5677), .C0(n6430), 
        .C1(n6503), .Y(n3693) );
  OAI222XL U8483 ( .A0(n6354), .A1(n5909), .B0(n3650), .B1(n3651), .C0(n638), 
        .C1(n3652), .Y(n4536) );
  AOI211X1 U8484 ( .A0(n5948), .A1(n3653), .B0(n3654), .C0(n5758), .Y(n3650)
         );
  OAI222XL U8485 ( .A0(n3655), .A1(n5702), .B0(n3656), .B1(n5677), .C0(n6431), 
        .C1(n5727), .Y(n3654) );
  OAI222XL U8486 ( .A0(n6355), .A1(n5909), .B0(n3611), .B1(n3612), .C0(n630), 
        .C1(n3613), .Y(n4528) );
  AOI211X1 U8487 ( .A0(n5948), .A1(n3614), .B0(n3615), .C0(n5760), .Y(n3611)
         );
  OAI222XL U8488 ( .A0(n3616), .A1(n5703), .B0(n3617), .B1(n5677), .C0(n6432), 
        .C1(n5729), .Y(n3615) );
  OAI222XL U8489 ( .A0(n6356), .A1(n5909), .B0(n3572), .B1(n3573), .C0(n622), 
        .C1(n3574), .Y(n4520) );
  AOI211X1 U8490 ( .A0(n5948), .A1(n3575), .B0(n3576), .C0(n5760), .Y(n3572)
         );
  OAI222XL U8491 ( .A0(n3577), .A1(n5702), .B0(n3578), .B1(n5677), .C0(n6433), 
        .C1(n5728), .Y(n3576) );
  OAI222XL U8492 ( .A0(n6357), .A1(n5909), .B0(n3533), .B1(n3534), .C0(n614), 
        .C1(n3535), .Y(n4512) );
  AOI211X1 U8493 ( .A0(n5948), .A1(n3536), .B0(n3537), .C0(n5760), .Y(n3533)
         );
  OAI222XL U8494 ( .A0(n3538), .A1(n5703), .B0(n3539), .B1(n5677), .C0(n6434), 
        .C1(n5727), .Y(n3537) );
  OAI222XL U8495 ( .A0(n6358), .A1(n5911), .B0(n3494), .B1(n3495), .C0(n606), 
        .C1(n3496), .Y(n4504) );
  AOI211X1 U8496 ( .A0(n5948), .A1(n3497), .B0(n3498), .C0(n5760), .Y(n3494)
         );
  OAI222XL U8497 ( .A0(n3499), .A1(n5702), .B0(n3500), .B1(n5677), .C0(n6435), 
        .C1(n5727), .Y(n3498) );
  OAI222XL U8498 ( .A0(n6359), .A1(n5910), .B0(n3455), .B1(n3456), .C0(n598), 
        .C1(n3457), .Y(n4496) );
  AOI211X1 U8499 ( .A0(n5948), .A1(n3458), .B0(n3459), .C0(n5760), .Y(n3455)
         );
  OAI222XL U8500 ( .A0(n3460), .A1(n5702), .B0(n3461), .B1(n5677), .C0(n6436), 
        .C1(n5727), .Y(n3459) );
  OAI222XL U8501 ( .A0(n6360), .A1(n5909), .B0(n3416), .B1(n3417), .C0(n590), 
        .C1(n3418), .Y(n4488) );
  AOI211X1 U8502 ( .A0(n5948), .A1(n3419), .B0(n3420), .C0(n5760), .Y(n3416)
         );
  OAI222XL U8503 ( .A0(n3421), .A1(n5702), .B0(n3422), .B1(n5677), .C0(n6437), 
        .C1(n5727), .Y(n3420) );
  OAI222XL U8504 ( .A0(n6361), .A1(n5911), .B0(n3372), .B1(n3373), .C0(n582), 
        .C1(n3374), .Y(n4480) );
  AOI211X1 U8505 ( .A0(n5948), .A1(n3375), .B0(n3376), .C0(n5760), .Y(n3372)
         );
  OAI222XL U8506 ( .A0(n3377), .A1(n5702), .B0(n3378), .B1(n5677), .C0(n6438), 
        .C1(n6503), .Y(n3376) );
  OAI222XL U8507 ( .A0(n6362), .A1(n5910), .B0(n3333), .B1(n3334), .C0(n574), 
        .C1(n3335), .Y(n4472) );
  AOI211X1 U8508 ( .A0(n5948), .A1(n3336), .B0(n3337), .C0(n5760), .Y(n3333)
         );
  OAI222XL U8509 ( .A0(n3338), .A1(n5702), .B0(n3339), .B1(n5677), .C0(n6439), 
        .C1(n5727), .Y(n3337) );
  OAI222XL U8510 ( .A0(n6363), .A1(n5909), .B0(n3294), .B1(n3295), .C0(n566), 
        .C1(n3296), .Y(n4464) );
  AOI211X1 U8511 ( .A0(n5948), .A1(n3297), .B0(n3298), .C0(n5760), .Y(n3294)
         );
  OAI222XL U8512 ( .A0(n3299), .A1(n5702), .B0(n3300), .B1(n5677), .C0(n6440), 
        .C1(n5727), .Y(n3298) );
  OAI222XL U8513 ( .A0(n6364), .A1(n5911), .B0(n3255), .B1(n3256), .C0(n558), 
        .C1(n3257), .Y(n4456) );
  AOI211X1 U8514 ( .A0(n5948), .A1(n3258), .B0(n3259), .C0(n5760), .Y(n3255)
         );
  OAI222XL U8515 ( .A0(n3260), .A1(n5702), .B0(n3261), .B1(n5675), .C0(n6441), 
        .C1(n6195), .Y(n3259) );
  OAI222XL U8516 ( .A0(n6365), .A1(n5910), .B0(n3216), .B1(n3217), .C0(n550), 
        .C1(n3218), .Y(n4448) );
  AOI211X1 U8517 ( .A0(n5948), .A1(n3219), .B0(n3220), .C0(n5760), .Y(n3216)
         );
  OAI222XL U8518 ( .A0(n3221), .A1(n5702), .B0(n3222), .B1(n5676), .C0(n6442), 
        .C1(n5729), .Y(n3220) );
  OAI222XL U8519 ( .A0(n6366), .A1(n5909), .B0(n3177), .B1(n3178), .C0(n542), 
        .C1(n3179), .Y(n4440) );
  AOI211X1 U8520 ( .A0(n5948), .A1(n3180), .B0(n3181), .C0(n5760), .Y(n3177)
         );
  OAI222XL U8521 ( .A0(n3182), .A1(n5702), .B0(n3183), .B1(n5675), .C0(n6443), 
        .C1(n5729), .Y(n3181) );
  OAI222XL U8522 ( .A0(n6367), .A1(n5909), .B0(n3138), .B1(n3139), .C0(n534), 
        .C1(n4674), .Y(n4432) );
  AOI211X1 U8523 ( .A0(n5948), .A1(n3141), .B0(n3142), .C0(n5760), .Y(n3138)
         );
  OAI222XL U8524 ( .A0(n3143), .A1(n5702), .B0(n3144), .B1(n5677), .C0(n6444), 
        .C1(n5729), .Y(n3142) );
  OAI222XL U8525 ( .A0(n6368), .A1(n5911), .B0(n3099), .B1(n3100), .C0(n526), 
        .C1(n3101), .Y(n4424) );
  AOI211X1 U8526 ( .A0(n5948), .A1(n3102), .B0(n3103), .C0(n5760), .Y(n3099)
         );
  OAI222XL U8527 ( .A0(n3104), .A1(n5702), .B0(n3105), .B1(n5675), .C0(n6445), 
        .C1(n5729), .Y(n3103) );
  OAI222XL U8528 ( .A0(n6369), .A1(n5910), .B0(n3055), .B1(n3056), .C0(n518), 
        .C1(n3057), .Y(n4416) );
  AOI211X1 U8529 ( .A0(n5948), .A1(n3058), .B0(n3059), .C0(n5760), .Y(n3055)
         );
  OAI222XL U8530 ( .A0(n3060), .A1(n5702), .B0(n3061), .B1(n5677), .C0(n6446), 
        .C1(n5729), .Y(n3059) );
  OAI222XL U8531 ( .A0(n6370), .A1(n5910), .B0(n3016), .B1(n3017), .C0(n510), 
        .C1(n3018), .Y(n4408) );
  AOI211X1 U8532 ( .A0(n5948), .A1(n3019), .B0(n3020), .C0(n5759), .Y(n3016)
         );
  OAI222XL U8533 ( .A0(n3021), .A1(n5704), .B0(n3022), .B1(n5675), .C0(n6447), 
        .C1(n5729), .Y(n3020) );
  OAI222XL U8534 ( .A0(n6371), .A1(n5910), .B0(n2977), .B1(n2978), .C0(n502), 
        .C1(n2979), .Y(n4400) );
  AOI211X1 U8535 ( .A0(n5948), .A1(n2980), .B0(n2981), .C0(n5759), .Y(n2977)
         );
  OAI222XL U8536 ( .A0(n2982), .A1(n5704), .B0(n2983), .B1(n5677), .C0(n6448), 
        .C1(n5729), .Y(n2981) );
  OAI222XL U8537 ( .A0(n6372), .A1(n5910), .B0(n2938), .B1(n2939), .C0(n494), 
        .C1(n4675), .Y(n4392) );
  AOI211X1 U8538 ( .A0(n5948), .A1(n2941), .B0(n2942), .C0(n5759), .Y(n2938)
         );
  OAI222XL U8539 ( .A0(n2943), .A1(n5704), .B0(n2944), .B1(n5676), .C0(n6449), 
        .C1(n5729), .Y(n2942) );
  OAI222XL U8540 ( .A0(n6373), .A1(n5910), .B0(n2899), .B1(n2900), .C0(n486), 
        .C1(n2901), .Y(n4384) );
  AOI211X1 U8541 ( .A0(n5948), .A1(n2902), .B0(n2903), .C0(n5759), .Y(n2899)
         );
  OAI222XL U8542 ( .A0(n2904), .A1(n5703), .B0(n2905), .B1(n5675), .C0(n6450), 
        .C1(n5729), .Y(n2903) );
  OAI222XL U8543 ( .A0(n6374), .A1(n5910), .B0(n2860), .B1(n2861), .C0(n478), 
        .C1(n2862), .Y(n4376) );
  AOI211X1 U8544 ( .A0(n5948), .A1(n2863), .B0(n2864), .C0(n5759), .Y(n2860)
         );
  OAI222XL U8545 ( .A0(n2865), .A1(n5704), .B0(n2866), .B1(n5677), .C0(n6451), 
        .C1(n5729), .Y(n2864) );
  OAI222XL U8546 ( .A0(n6375), .A1(n5910), .B0(n2821), .B1(n2822), .C0(n470), 
        .C1(n2823), .Y(n4368) );
  AOI211X1 U8547 ( .A0(n5948), .A1(n2824), .B0(n2825), .C0(n5759), .Y(n2821)
         );
  OAI222XL U8548 ( .A0(n2826), .A1(n5703), .B0(n2827), .B1(n6007), .C0(n6452), 
        .C1(n5729), .Y(n2825) );
  OAI222XL U8549 ( .A0(n6376), .A1(n5910), .B0(n2782), .B1(n2783), .C0(n462), 
        .C1(n2784), .Y(n4360) );
  AOI211X1 U8550 ( .A0(n5948), .A1(n2785), .B0(n2786), .C0(n5759), .Y(n2782)
         );
  OAI222XL U8551 ( .A0(n2787), .A1(n5704), .B0(n2788), .B1(n6007), .C0(n6453), 
        .C1(n5729), .Y(n2786) );
  OAI222XL U8552 ( .A0(n6377), .A1(n5910), .B0(n2738), .B1(n2739), .C0(n454), 
        .C1(n2740), .Y(n4352) );
  AOI211X1 U8553 ( .A0(n5948), .A1(n2741), .B0(n2742), .C0(n5759), .Y(n2738)
         );
  OAI222XL U8554 ( .A0(n2743), .A1(n5704), .B0(n2744), .B1(n5677), .C0(n6454), 
        .C1(n5729), .Y(n2742) );
  OAI222XL U8555 ( .A0(n6378), .A1(n5910), .B0(n2699), .B1(n2700), .C0(n446), 
        .C1(n2701), .Y(n4344) );
  AOI211X1 U8556 ( .A0(n5948), .A1(n2702), .B0(n2703), .C0(n5759), .Y(n2699)
         );
  OAI222XL U8557 ( .A0(n2704), .A1(n5703), .B0(n2705), .B1(n6007), .C0(n6455), 
        .C1(n5729), .Y(n2703) );
  OAI222XL U8558 ( .A0(n6379), .A1(n5910), .B0(n2660), .B1(n2661), .C0(n438), 
        .C1(n2662), .Y(n4336) );
  AOI211X1 U8559 ( .A0(n5948), .A1(n2663), .B0(n2664), .C0(n5759), .Y(n2660)
         );
  OAI222XL U8560 ( .A0(n2665), .A1(n5704), .B0(n2666), .B1(n5676), .C0(n6456), 
        .C1(n5729), .Y(n2664) );
  OAI222XL U8561 ( .A0(n6380), .A1(n5910), .B0(n2621), .B1(n2622), .C0(n430), 
        .C1(n2623), .Y(n4328) );
  AOI211X1 U8562 ( .A0(n5948), .A1(n2624), .B0(n2625), .C0(n5759), .Y(n2621)
         );
  OAI222XL U8563 ( .A0(n2626), .A1(n5703), .B0(n2627), .B1(n5676), .C0(n6457), 
        .C1(n6228), .Y(n2625) );
  OAI222XL U8564 ( .A0(n6381), .A1(n5910), .B0(n2582), .B1(n2583), .C0(n422), 
        .C1(n2584), .Y(n4320) );
  AOI211X1 U8565 ( .A0(n5948), .A1(n2585), .B0(n2586), .C0(n5759), .Y(n2582)
         );
  OAI222XL U8566 ( .A0(n2587), .A1(n5702), .B0(n2588), .B1(n5676), .C0(n6458), 
        .C1(n6228), .Y(n2586) );
  OAI222XL U8567 ( .A0(n6382), .A1(n5911), .B0(n2543), .B1(n2544), .C0(n414), 
        .C1(n2545), .Y(n4312) );
  AOI211X1 U8568 ( .A0(n5948), .A1(n2546), .B0(n2547), .C0(n5759), .Y(n2543)
         );
  OAI222XL U8569 ( .A0(n2548), .A1(n5703), .B0(n2549), .B1(n5676), .C0(n6459), 
        .C1(n6260), .Y(n2547) );
  OAI222XL U8570 ( .A0(n6383), .A1(n5911), .B0(n2504), .B1(n2505), .C0(n406), 
        .C1(n2506), .Y(n4304) );
  AOI211X1 U8571 ( .A0(n5948), .A1(n2507), .B0(n2508), .C0(n5758), .Y(n2504)
         );
  OAI222XL U8572 ( .A0(n2509), .A1(n5703), .B0(n2510), .B1(n5676), .C0(n6460), 
        .C1(n6195), .Y(n2508) );
  OAI222XL U8573 ( .A0(n6384), .A1(n5911), .B0(n2465), .B1(n2466), .C0(n398), 
        .C1(n2467), .Y(n4296) );
  AOI211X1 U8574 ( .A0(n5948), .A1(n2468), .B0(n2469), .C0(n5758), .Y(n2465)
         );
  OAI222XL U8575 ( .A0(n2470), .A1(n5703), .B0(n2471), .B1(n5676), .C0(n6461), 
        .C1(n5728), .Y(n2469) );
  OAI222XL U8576 ( .A0(n6385), .A1(n5911), .B0(n2421), .B1(n2422), .C0(n390), 
        .C1(n2423), .Y(n4288) );
  AOI211X1 U8577 ( .A0(n5948), .A1(n2424), .B0(n2425), .C0(n5758), .Y(n2421)
         );
  OAI222XL U8578 ( .A0(n2426), .A1(n5703), .B0(n2427), .B1(n5676), .C0(n6462), 
        .C1(n5727), .Y(n2425) );
  OAI222XL U8579 ( .A0(n6386), .A1(n5911), .B0(n2382), .B1(n2383), .C0(n382), 
        .C1(n2384), .Y(n4280) );
  AOI211X1 U8580 ( .A0(n5948), .A1(n2385), .B0(n2386), .C0(n5758), .Y(n2382)
         );
  OAI222XL U8581 ( .A0(n2387), .A1(n5703), .B0(n2388), .B1(n5676), .C0(n6463), 
        .C1(n6260), .Y(n2386) );
  OAI222XL U8582 ( .A0(n6387), .A1(n5911), .B0(n2343), .B1(n2344), .C0(n374), 
        .C1(n2345), .Y(n4272) );
  AOI211X1 U8583 ( .A0(n5948), .A1(n2346), .B0(n2347), .C0(n5758), .Y(n2343)
         );
  OAI222XL U8584 ( .A0(n2348), .A1(n5703), .B0(n2349), .B1(n5676), .C0(n6464), 
        .C1(n5727), .Y(n2347) );
  OAI222XL U8585 ( .A0(n6388), .A1(n5911), .B0(n2304), .B1(n2305), .C0(n366), 
        .C1(n2306), .Y(n4264) );
  AOI211X1 U8586 ( .A0(n5948), .A1(n2307), .B0(n2308), .C0(n5758), .Y(n2304)
         );
  OAI222XL U8587 ( .A0(n2309), .A1(n5703), .B0(n2310), .B1(n5676), .C0(n6465), 
        .C1(n6228), .Y(n2308) );
  OAI222XL U8588 ( .A0(n6389), .A1(n5911), .B0(n2265), .B1(n2266), .C0(n358), 
        .C1(n2267), .Y(n4256) );
  AOI211X1 U8589 ( .A0(n5948), .A1(n2268), .B0(n2269), .C0(n5758), .Y(n2265)
         );
  OAI222XL U8590 ( .A0(n2270), .A1(n5703), .B0(n2271), .B1(n5676), .C0(n6466), 
        .C1(n6195), .Y(n2269) );
  OAI222XL U8591 ( .A0(n6390), .A1(n5911), .B0(n2226), .B1(n2227), .C0(n350), 
        .C1(n2228), .Y(n4248) );
  AOI211X1 U8592 ( .A0(n5948), .A1(n2229), .B0(n2230), .C0(n5758), .Y(n2226)
         );
  OAI222XL U8593 ( .A0(n2231), .A1(n5703), .B0(n2232), .B1(n5676), .C0(n6467), 
        .C1(n5727), .Y(n2230) );
  OAI222XL U8594 ( .A0(n6391), .A1(n5911), .B0(n2187), .B1(n2188), .C0(n342), 
        .C1(n2189), .Y(n4240) );
  AOI211X1 U8595 ( .A0(n5948), .A1(n2190), .B0(n2191), .C0(n5758), .Y(n2187)
         );
  OAI222XL U8596 ( .A0(n2192), .A1(n5703), .B0(n2193), .B1(n5676), .C0(n6468), 
        .C1(n6260), .Y(n2191) );
  OAI222XL U8597 ( .A0(n6392), .A1(n5911), .B0(n2148), .B1(n2149), .C0(n334), 
        .C1(n2150), .Y(n4232) );
  AOI211X1 U8598 ( .A0(n5948), .A1(n2151), .B0(n2152), .C0(n5758), .Y(n2148)
         );
  OAI222XL U8599 ( .A0(n2153), .A1(n5703), .B0(n2154), .B1(n5676), .C0(n6469), 
        .C1(n5729), .Y(n2152) );
  OAI222XL U8600 ( .A0(n6393), .A1(n5911), .B0(n2104), .B1(n2105), .C0(n326), 
        .C1(n2106), .Y(n4224) );
  AOI211X1 U8601 ( .A0(n5948), .A1(n2107), .B0(n2108), .C0(n5758), .Y(n2104)
         );
  OAI222XL U8602 ( .A0(n2109), .A1(n5703), .B0(n2110), .B1(n5676), .C0(n6470), 
        .C1(n5729), .Y(n2108) );
  OAI222XL U8603 ( .A0(n6394), .A1(n5909), .B0(n2065), .B1(n2066), .C0(n318), 
        .C1(n2067), .Y(n4216) );
  AOI211X1 U8604 ( .A0(n5948), .A1(n2068), .B0(n2069), .C0(n5758), .Y(n2065)
         );
  OAI222XL U8605 ( .A0(n2070), .A1(n5704), .B0(n2071), .B1(n5676), .C0(n6471), 
        .C1(n6503), .Y(n2069) );
  OAI222XL U8606 ( .A0(n6395), .A1(n5909), .B0(n2026), .B1(n2027), .C0(n310), 
        .C1(n2028), .Y(n4208) );
  AOI211X1 U8607 ( .A0(n5948), .A1(n2029), .B0(n2030), .C0(n5758), .Y(n2026)
         );
  OAI222XL U8608 ( .A0(n2031), .A1(n5704), .B0(n2032), .B1(n5675), .C0(n6472), 
        .C1(n6228), .Y(n2030) );
  OAI222XL U8609 ( .A0(n6396), .A1(n5911), .B0(n1986), .B1(n1987), .C0(n302), 
        .C1(n1988), .Y(n4200) );
  AOI211X1 U8610 ( .A0(n5948), .A1(n6473), .B0(n1989), .C0(n5759), .Y(n1986)
         );
  OAI222XL U8611 ( .A0(n1990), .A1(n5704), .B0(n1991), .B1(n5675), .C0(n6474), 
        .C1(n5728), .Y(n1989) );
  OAI222XL U8612 ( .A0(n6397), .A1(n5911), .B0(n1947), .B1(n1948), .C0(n294), 
        .C1(n1949), .Y(n4192) );
  AOI211X1 U8613 ( .A0(n5948), .A1(n6475), .B0(n1950), .C0(n5758), .Y(n1947)
         );
  OAI222XL U8614 ( .A0(n1951), .A1(n5704), .B0(n1952), .B1(n5675), .C0(n6476), 
        .C1(n5728), .Y(n1950) );
  OAI222XL U8615 ( .A0(n6398), .A1(n5911), .B0(n1908), .B1(n1909), .C0(n286), 
        .C1(n1910), .Y(n4184) );
  AOI211X1 U8616 ( .A0(n5948), .A1(n6477), .B0(n1911), .C0(n5760), .Y(n1908)
         );
  OAI222XL U8617 ( .A0(n1912), .A1(n5704), .B0(n1913), .B1(n5675), .C0(n6478), 
        .C1(n5728), .Y(n1911) );
  OAI222XL U8618 ( .A0(n4832), .A1(n5910), .B0(n1869), .B1(n1870), .C0(n278), 
        .C1(n1871), .Y(n4176) );
  AOI211X1 U8619 ( .A0(n5948), .A1(n6479), .B0(n1872), .C0(n5759), .Y(n1869)
         );
  OAI222XL U8620 ( .A0(n1873), .A1(n5704), .B0(n1874), .B1(n5675), .C0(n6480), 
        .C1(n5728), .Y(n1872) );
  OAI222XL U8621 ( .A0(n6399), .A1(n5910), .B0(n1830), .B1(n1831), .C0(n270), 
        .C1(n4643), .Y(n4168) );
  AOI211X1 U8622 ( .A0(n5948), .A1(n6481), .B0(n1833), .C0(n5758), .Y(n1830)
         );
  OAI222XL U8623 ( .A0(n1834), .A1(n5704), .B0(n1835), .B1(n5675), .C0(n6482), 
        .C1(n5728), .Y(n1833) );
  OAI222XL U8624 ( .A0(n6400), .A1(n5910), .B0(n1786), .B1(n1787), .C0(n262), 
        .C1(n1788), .Y(n4160) );
  AOI211X1 U8625 ( .A0(n5948), .A1(n6483), .B0(n1789), .C0(n5760), .Y(n1786)
         );
  OAI222XL U8626 ( .A0(n1790), .A1(n5704), .B0(n1791), .B1(n5675), .C0(n6484), 
        .C1(n5728), .Y(n1789) );
  OAI222XL U8627 ( .A0(n6401), .A1(n5909), .B0(n1741), .B1(n1742), .C0(n254), 
        .C1(n1743), .Y(n4152) );
  AOI211X1 U8628 ( .A0(n5948), .A1(n6485), .B0(n1744), .C0(n5759), .Y(n1741)
         );
  OAI222XL U8629 ( .A0(n1745), .A1(n5704), .B0(n1746), .B1(n5675), .C0(n6486), 
        .C1(n5728), .Y(n1744) );
  OAI222XL U8630 ( .A0(n6402), .A1(n5911), .B0(n1697), .B1(n1698), .C0(n246), 
        .C1(n1699), .Y(n4144) );
  AOI211X1 U8631 ( .A0(n5948), .A1(n6487), .B0(n1700), .C0(n5758), .Y(n1697)
         );
  OAI222XL U8632 ( .A0(n1701), .A1(n5704), .B0(n1702), .B1(n5675), .C0(n6488), 
        .C1(n5728), .Y(n1700) );
  OAI222XL U8633 ( .A0(n6403), .A1(n5910), .B0(n1653), .B1(n1654), .C0(n238), 
        .C1(n1655), .Y(n4136) );
  AOI211X1 U8634 ( .A0(n5948), .A1(n6489), .B0(n1656), .C0(n5760), .Y(n1653)
         );
  OAI222XL U8635 ( .A0(n1657), .A1(n5704), .B0(n1658), .B1(n5675), .C0(n6490), 
        .C1(n5728), .Y(n1656) );
  OAI222XL U8636 ( .A0(n6404), .A1(n5910), .B0(n1609), .B1(n1610), .C0(n230), 
        .C1(n1611), .Y(n4128) );
  AOI211X1 U8637 ( .A0(n5948), .A1(n6491), .B0(n1612), .C0(n5759), .Y(n1609)
         );
  OAI222XL U8638 ( .A0(n1613), .A1(n5704), .B0(n1614), .B1(n5675), .C0(n6492), 
        .C1(n5728), .Y(n1612) );
  OAI222XL U8639 ( .A0(n6405), .A1(n5909), .B0(n1565), .B1(n1566), .C0(n222), 
        .C1(n1567), .Y(n4120) );
  AOI211X1 U8640 ( .A0(n5948), .A1(n6493), .B0(n1568), .C0(n5758), .Y(n1565)
         );
  OAI222XL U8641 ( .A0(n1569), .A1(n5702), .B0(n1570), .B1(n5675), .C0(n6494), 
        .C1(n5728), .Y(n1568) );
  OAI222XL U8642 ( .A0(n6406), .A1(n5909), .B0(n1521), .B1(n1522), .C0(n214), 
        .C1(n1523), .Y(n4112) );
  AOI211X1 U8643 ( .A0(n5948), .A1(n6495), .B0(n1524), .C0(n5760), .Y(n1521)
         );
  OAI222XL U8644 ( .A0(n1525), .A1(n5702), .B0(n1526), .B1(n5675), .C0(n6496), 
        .C1(n5728), .Y(n1524) );
  OAI222XL U8645 ( .A0(n6407), .A1(n5911), .B0(n1477), .B1(n1478), .C0(n206), 
        .C1(n1479), .Y(n4104) );
  AOI211X1 U8646 ( .A0(n5948), .A1(n6497), .B0(n1480), .C0(n5759), .Y(n1477)
         );
  OAI222XL U8647 ( .A0(n1481), .A1(n5704), .B0(n1482), .B1(n5676), .C0(n6498), 
        .C1(n5729), .Y(n1480) );
  OAI222XL U8648 ( .A0(n6347), .A1(n5906), .B0(n3935), .B1(n3929), .C0(n695), 
        .C1(n3930), .Y(n4593) );
  AOI211X1 U8649 ( .A0(n5944), .A1(n3931), .B0(n3936), .C0(n5755), .Y(n3935)
         );
  OAI222XL U8650 ( .A0(n3933), .A1(n5705), .B0(n3934), .B1(n5678), .C0(n6424), 
        .C1(n5731), .Y(n3936) );
  OAI222XL U8651 ( .A0(n6348), .A1(n5906), .B0(n3896), .B1(n3890), .C0(n687), 
        .C1(n3891), .Y(n4585) );
  AOI211X1 U8652 ( .A0(n5944), .A1(n3892), .B0(n3897), .C0(n5755), .Y(n3896)
         );
  OAI222XL U8653 ( .A0(n3894), .A1(n5705), .B0(n3895), .B1(n5680), .C0(n6425), 
        .C1(n5731), .Y(n3897) );
  OAI222XL U8654 ( .A0(n6349), .A1(n5906), .B0(n3857), .B1(n3851), .C0(n679), 
        .C1(n3852), .Y(n4577) );
  AOI211X1 U8655 ( .A0(n5944), .A1(n3853), .B0(n3858), .C0(n5755), .Y(n3857)
         );
  OAI222XL U8656 ( .A0(n3855), .A1(n5705), .B0(n3856), .B1(n5680), .C0(n6426), 
        .C1(n5732), .Y(n3858) );
  OAI222XL U8657 ( .A0(n6350), .A1(n5906), .B0(n3818), .B1(n3812), .C0(n671), 
        .C1(n3813), .Y(n4569) );
  AOI211X1 U8658 ( .A0(n5944), .A1(n3814), .B0(n3819), .C0(n5755), .Y(n3818)
         );
  OAI222XL U8659 ( .A0(n3816), .A1(n5705), .B0(n3817), .B1(n5680), .C0(n6427), 
        .C1(n5732), .Y(n3819) );
  OAI222XL U8660 ( .A0(n6351), .A1(n5906), .B0(n3779), .B1(n3773), .C0(n663), 
        .C1(n3774), .Y(n4561) );
  AOI211X1 U8661 ( .A0(n5944), .A1(n3775), .B0(n3780), .C0(n5755), .Y(n3779)
         );
  OAI222XL U8662 ( .A0(n3777), .A1(n5705), .B0(n3778), .B1(n5680), .C0(n6428), 
        .C1(n5732), .Y(n3780) );
  OAI222XL U8663 ( .A0(n6352), .A1(n5906), .B0(n3740), .B1(n3734), .C0(n655), 
        .C1(n3735), .Y(n4553) );
  AOI211X1 U8664 ( .A0(n5944), .A1(n3736), .B0(n3741), .C0(n5755), .Y(n3740)
         );
  OAI222XL U8665 ( .A0(n3738), .A1(n5705), .B0(n3739), .B1(n5680), .C0(n6429), 
        .C1(n5732), .Y(n3741) );
  OAI222XL U8666 ( .A0(n6353), .A1(n5906), .B0(n3696), .B1(n3690), .C0(n647), 
        .C1(n5670), .Y(n4545) );
  AOI211X1 U8667 ( .A0(n5944), .A1(n3692), .B0(n3697), .C0(n5755), .Y(n3696)
         );
  OAI222XL U8668 ( .A0(n3694), .A1(n5705), .B0(n3695), .B1(n5680), .C0(n6430), 
        .C1(n5730), .Y(n3697) );
  OAI222XL U8669 ( .A0(n6354), .A1(n5906), .B0(n3657), .B1(n3651), .C0(n639), 
        .C1(n3652), .Y(n4537) );
  AOI211X1 U8670 ( .A0(n5944), .A1(n3653), .B0(n3658), .C0(n5755), .Y(n3657)
         );
  OAI222XL U8671 ( .A0(n3655), .A1(n5705), .B0(n3656), .B1(n5680), .C0(n6431), 
        .C1(n5730), .Y(n3658) );
  OAI222XL U8672 ( .A0(n6355), .A1(n5906), .B0(n3618), .B1(n3612), .C0(n631), 
        .C1(n3613), .Y(n4529) );
  AOI211X1 U8673 ( .A0(n5944), .A1(n3614), .B0(n3619), .C0(n5755), .Y(n3618)
         );
  OAI222XL U8674 ( .A0(n3616), .A1(n5705), .B0(n3617), .B1(n5680), .C0(n6432), 
        .C1(n5731), .Y(n3619) );
  OAI222XL U8675 ( .A0(n6356), .A1(n5906), .B0(n3579), .B1(n3573), .C0(n623), 
        .C1(n3574), .Y(n4521) );
  AOI211X1 U8676 ( .A0(n5944), .A1(n3575), .B0(n3580), .C0(n5755), .Y(n3579)
         );
  OAI222XL U8677 ( .A0(n3577), .A1(n5705), .B0(n3578), .B1(n5680), .C0(n6433), 
        .C1(n5731), .Y(n3580) );
  OAI222XL U8678 ( .A0(n6357), .A1(n5906), .B0(n3540), .B1(n3534), .C0(n615), 
        .C1(n3535), .Y(n4513) );
  AOI211X1 U8679 ( .A0(n5944), .A1(n3536), .B0(n3541), .C0(n5754), .Y(n3540)
         );
  OAI222XL U8680 ( .A0(n3538), .A1(n5705), .B0(n3539), .B1(n5680), .C0(n6434), 
        .C1(n5732), .Y(n3541) );
  OAI222XL U8681 ( .A0(n6358), .A1(n5906), .B0(n3501), .B1(n3495), .C0(n607), 
        .C1(n3496), .Y(n4505) );
  AOI211X1 U8682 ( .A0(n5944), .A1(n3497), .B0(n3502), .C0(n5754), .Y(n3501)
         );
  OAI222XL U8683 ( .A0(n3499), .A1(n5706), .B0(n3500), .B1(n5680), .C0(n6435), 
        .C1(n5731), .Y(n3502) );
  OAI222XL U8684 ( .A0(n6359), .A1(n5907), .B0(n3462), .B1(n3456), .C0(n599), 
        .C1(n3457), .Y(n4497) );
  AOI211X1 U8685 ( .A0(n5944), .A1(n3458), .B0(n3463), .C0(n5754), .Y(n3462)
         );
  OAI222XL U8686 ( .A0(n3460), .A1(n5706), .B0(n3461), .B1(n5680), .C0(n6436), 
        .C1(n6504), .Y(n3463) );
  OAI222XL U8687 ( .A0(n6360), .A1(n5908), .B0(n3423), .B1(n3417), .C0(n591), 
        .C1(n3418), .Y(n4489) );
  AOI211X1 U8688 ( .A0(n5944), .A1(n3419), .B0(n3424), .C0(n5754), .Y(n3423)
         );
  OAI222XL U8689 ( .A0(n3421), .A1(n5706), .B0(n3422), .B1(n5680), .C0(n6437), 
        .C1(n6504), .Y(n3424) );
  OAI222XL U8690 ( .A0(n6361), .A1(n5906), .B0(n3379), .B1(n3373), .C0(n583), 
        .C1(n3374), .Y(n4481) );
  AOI211X1 U8691 ( .A0(n5944), .A1(n3375), .B0(n3380), .C0(n5754), .Y(n3379)
         );
  OAI222XL U8692 ( .A0(n3377), .A1(n5706), .B0(n3378), .B1(n5680), .C0(n6438), 
        .C1(n6504), .Y(n3380) );
  OAI222XL U8693 ( .A0(n6362), .A1(n5907), .B0(n3340), .B1(n3334), .C0(n575), 
        .C1(n3335), .Y(n4473) );
  AOI211X1 U8694 ( .A0(n5944), .A1(n3336), .B0(n3341), .C0(n5754), .Y(n3340)
         );
  OAI222XL U8695 ( .A0(n3338), .A1(n5706), .B0(n3339), .B1(n5680), .C0(n6439), 
        .C1(n6504), .Y(n3341) );
  OAI222XL U8696 ( .A0(n6363), .A1(n5908), .B0(n3301), .B1(n3295), .C0(n567), 
        .C1(n3296), .Y(n4465) );
  AOI211X1 U8697 ( .A0(n5944), .A1(n3297), .B0(n3302), .C0(n5754), .Y(n3301)
         );
  OAI222XL U8698 ( .A0(n3299), .A1(n5706), .B0(n3300), .B1(n5680), .C0(n6440), 
        .C1(n6504), .Y(n3302) );
  OAI222XL U8699 ( .A0(n6364), .A1(n5906), .B0(n3262), .B1(n3256), .C0(n559), 
        .C1(n3257), .Y(n4457) );
  AOI211X1 U8700 ( .A0(n5944), .A1(n3258), .B0(n3263), .C0(n5754), .Y(n3262)
         );
  OAI222XL U8701 ( .A0(n3260), .A1(n5706), .B0(n3261), .B1(n5680), .C0(n6441), 
        .C1(n6504), .Y(n3263) );
  OAI222XL U8702 ( .A0(n6365), .A1(n5907), .B0(n3223), .B1(n3217), .C0(n551), 
        .C1(n3218), .Y(n4449) );
  AOI211X1 U8703 ( .A0(n5944), .A1(n3219), .B0(n3224), .C0(n5754), .Y(n3223)
         );
  OAI222XL U8704 ( .A0(n3221), .A1(n5706), .B0(n3222), .B1(n5680), .C0(n6442), 
        .C1(n5732), .Y(n3224) );
  OAI222XL U8705 ( .A0(n6366), .A1(n5908), .B0(n3184), .B1(n3178), .C0(n543), 
        .C1(n3179), .Y(n4441) );
  AOI211X1 U8706 ( .A0(n5944), .A1(n3180), .B0(n3185), .C0(n5754), .Y(n3184)
         );
  OAI222XL U8707 ( .A0(n3182), .A1(n5706), .B0(n3183), .B1(n5680), .C0(n6443), 
        .C1(n5732), .Y(n3185) );
  OAI222XL U8708 ( .A0(n6367), .A1(n5908), .B0(n3145), .B1(n3139), .C0(n535), 
        .C1(n4674), .Y(n4433) );
  AOI211X1 U8709 ( .A0(n5944), .A1(n3141), .B0(n3146), .C0(n5754), .Y(n3145)
         );
  OAI222XL U8710 ( .A0(n3143), .A1(n5706), .B0(n3144), .B1(n5678), .C0(n6444), 
        .C1(n5732), .Y(n3146) );
  OAI222XL U8711 ( .A0(n6368), .A1(n5906), .B0(n3106), .B1(n3100), .C0(n527), 
        .C1(n3101), .Y(n4425) );
  AOI211X1 U8712 ( .A0(n5944), .A1(n3102), .B0(n3107), .C0(n5754), .Y(n3106)
         );
  OAI222XL U8713 ( .A0(n3104), .A1(n5706), .B0(n3105), .B1(n5680), .C0(n6445), 
        .C1(n5732), .Y(n3107) );
  OAI222XL U8714 ( .A0(n6369), .A1(n5907), .B0(n3062), .B1(n3056), .C0(n519), 
        .C1(n3057), .Y(n4417) );
  AOI211X1 U8715 ( .A0(n5944), .A1(n3058), .B0(n3063), .C0(n5754), .Y(n3062)
         );
  OAI222XL U8716 ( .A0(n3060), .A1(n5706), .B0(n3061), .B1(n5679), .C0(n6446), 
        .C1(n5732), .Y(n3063) );
  OAI222XL U8717 ( .A0(n6370), .A1(n5907), .B0(n3023), .B1(n3017), .C0(n511), 
        .C1(n3018), .Y(n4409) );
  AOI211X1 U8718 ( .A0(n5944), .A1(n3019), .B0(n3024), .C0(n5753), .Y(n3023)
         );
  OAI222XL U8719 ( .A0(n3021), .A1(n5707), .B0(n3022), .B1(n6068), .C0(n6447), 
        .C1(n5732), .Y(n3024) );
  OAI222XL U8720 ( .A0(n6371), .A1(n5907), .B0(n2984), .B1(n2978), .C0(n503), 
        .C1(n2979), .Y(n4401) );
  AOI211X1 U8721 ( .A0(n5944), .A1(n2980), .B0(n2985), .C0(n5753), .Y(n2984)
         );
  OAI222XL U8722 ( .A0(n2982), .A1(n5705), .B0(n2983), .B1(n5678), .C0(n6448), 
        .C1(n5732), .Y(n2985) );
  OAI222XL U8723 ( .A0(n6372), .A1(n5907), .B0(n2945), .B1(n2939), .C0(n495), 
        .C1(n4675), .Y(n4393) );
  AOI211X1 U8724 ( .A0(n5944), .A1(n2941), .B0(n2946), .C0(n5753), .Y(n2945)
         );
  OAI222XL U8725 ( .A0(n2943), .A1(n5705), .B0(n2944), .B1(n5678), .C0(n6449), 
        .C1(n5732), .Y(n2946) );
  OAI222XL U8726 ( .A0(n6373), .A1(n5907), .B0(n2906), .B1(n2900), .C0(n487), 
        .C1(n2901), .Y(n4385) );
  AOI211X1 U8727 ( .A0(n5944), .A1(n2902), .B0(n2907), .C0(n5753), .Y(n2906)
         );
  OAI222XL U8728 ( .A0(n2904), .A1(n5707), .B0(n2905), .B1(n6417), .C0(n6450), 
        .C1(n5732), .Y(n2907) );
  OAI222XL U8729 ( .A0(n6374), .A1(n5907), .B0(n2867), .B1(n2861), .C0(n479), 
        .C1(n2862), .Y(n4377) );
  AOI211X1 U8730 ( .A0(n5944), .A1(n2863), .B0(n2868), .C0(n5753), .Y(n2867)
         );
  OAI222XL U8731 ( .A0(n2865), .A1(n5705), .B0(n2866), .B1(n6417), .C0(n6451), 
        .C1(n5732), .Y(n2868) );
  OAI222XL U8732 ( .A0(n6375), .A1(n5907), .B0(n2828), .B1(n2822), .C0(n471), 
        .C1(n2823), .Y(n4369) );
  AOI211X1 U8733 ( .A0(n5944), .A1(n2824), .B0(n2829), .C0(n5753), .Y(n2828)
         );
  OAI222XL U8734 ( .A0(n2826), .A1(n5706), .B0(n2827), .B1(n6417), .C0(n6452), 
        .C1(n5732), .Y(n2829) );
  OAI222XL U8735 ( .A0(n6376), .A1(n5907), .B0(n2789), .B1(n2783), .C0(n463), 
        .C1(n2784), .Y(n4361) );
  AOI211X1 U8736 ( .A0(n5944), .A1(n2785), .B0(n2790), .C0(n5753), .Y(n2789)
         );
  OAI222XL U8737 ( .A0(n2787), .A1(n5707), .B0(n2788), .B1(n6417), .C0(n6453), 
        .C1(n5732), .Y(n2790) );
  OAI222XL U8738 ( .A0(n6377), .A1(n5907), .B0(n2745), .B1(n2739), .C0(n455), 
        .C1(n2740), .Y(n4353) );
  AOI211X1 U8739 ( .A0(n5945), .A1(n2741), .B0(n2746), .C0(n5753), .Y(n2745)
         );
  OAI222XL U8740 ( .A0(n2743), .A1(n5705), .B0(n2744), .B1(n5678), .C0(n6454), 
        .C1(n5732), .Y(n2746) );
  OAI222XL U8741 ( .A0(n6378), .A1(n5907), .B0(n2706), .B1(n2700), .C0(n447), 
        .C1(n2701), .Y(n4345) );
  AOI211X1 U8742 ( .A0(n5944), .A1(n2702), .B0(n2707), .C0(n5753), .Y(n2706)
         );
  OAI222XL U8743 ( .A0(n2704), .A1(n5705), .B0(n2705), .B1(n6417), .C0(n6455), 
        .C1(n5732), .Y(n2707) );
  OAI222XL U8744 ( .A0(n6379), .A1(n5907), .B0(n2667), .B1(n2661), .C0(n439), 
        .C1(n2662), .Y(n4337) );
  AOI211X1 U8745 ( .A0(n5944), .A1(n2663), .B0(n2668), .C0(n5753), .Y(n2667)
         );
  OAI222XL U8746 ( .A0(n2665), .A1(n5707), .B0(n2666), .B1(n5678), .C0(n6456), 
        .C1(n5732), .Y(n2668) );
  OAI222XL U8747 ( .A0(n6380), .A1(n5907), .B0(n2628), .B1(n2622), .C0(n431), 
        .C1(n2623), .Y(n4329) );
  AOI211X1 U8748 ( .A0(n5945), .A1(n2624), .B0(n2629), .C0(n5753), .Y(n2628)
         );
  OAI222XL U8749 ( .A0(n2626), .A1(n5705), .B0(n2627), .B1(n5678), .C0(n6457), 
        .C1(n5730), .Y(n2629) );
  OAI222XL U8750 ( .A0(n6381), .A1(n5907), .B0(n2589), .B1(n2583), .C0(n423), 
        .C1(n2584), .Y(n4321) );
  AOI211X1 U8751 ( .A0(n5945), .A1(n2585), .B0(n2590), .C0(n5753), .Y(n2589)
         );
  OAI222XL U8752 ( .A0(n2587), .A1(n5705), .B0(n2588), .B1(n5678), .C0(n6458), 
        .C1(n5731), .Y(n2590) );
  OAI222XL U8753 ( .A0(n6382), .A1(n5908), .B0(n2550), .B1(n2544), .C0(n415), 
        .C1(n2545), .Y(n4313) );
  AOI211X1 U8754 ( .A0(n5945), .A1(n2546), .B0(n2551), .C0(n5753), .Y(n2550)
         );
  OAI222XL U8755 ( .A0(n2548), .A1(n5707), .B0(n2549), .B1(n5678), .C0(n6459), 
        .C1(n5731), .Y(n2551) );
  OAI222XL U8756 ( .A0(n6383), .A1(n5908), .B0(n2511), .B1(n2505), .C0(n407), 
        .C1(n2506), .Y(n4305) );
  AOI211X1 U8757 ( .A0(n5945), .A1(n2507), .B0(n2512), .C0(n5752), .Y(n2511)
         );
  OAI222XL U8758 ( .A0(n2509), .A1(n5707), .B0(n2510), .B1(n6417), .C0(n6460), 
        .C1(n5731), .Y(n2512) );
  OAI222XL U8759 ( .A0(n6384), .A1(n5908), .B0(n2472), .B1(n2466), .C0(n399), 
        .C1(n2467), .Y(n4297) );
  AOI211X1 U8760 ( .A0(n5945), .A1(n2468), .B0(n2473), .C0(n5752), .Y(n2472)
         );
  OAI222XL U8761 ( .A0(n2470), .A1(n5707), .B0(n2471), .B1(n5678), .C0(n6461), 
        .C1(n5731), .Y(n2473) );
  OAI222XL U8762 ( .A0(n6385), .A1(n5908), .B0(n2428), .B1(n2422), .C0(n391), 
        .C1(n2423), .Y(n4289) );
  AOI211X1 U8763 ( .A0(n5945), .A1(n2424), .B0(n2429), .C0(n5752), .Y(n2428)
         );
  OAI222XL U8764 ( .A0(n2426), .A1(n5707), .B0(n2427), .B1(n5678), .C0(n6462), 
        .C1(n5731), .Y(n2429) );
  OAI222XL U8765 ( .A0(n6386), .A1(n5908), .B0(n2389), .B1(n2383), .C0(n383), 
        .C1(n2384), .Y(n4281) );
  AOI211X1 U8766 ( .A0(n5945), .A1(n2385), .B0(n2390), .C0(n5752), .Y(n2389)
         );
  OAI222XL U8767 ( .A0(n2387), .A1(n5707), .B0(n2388), .B1(n5678), .C0(n6463), 
        .C1(n5731), .Y(n2390) );
  OAI222XL U8768 ( .A0(n6387), .A1(n5908), .B0(n2350), .B1(n2344), .C0(n375), 
        .C1(n2345), .Y(n4273) );
  AOI211X1 U8769 ( .A0(n5945), .A1(n2346), .B0(n2351), .C0(n5752), .Y(n2350)
         );
  OAI222XL U8770 ( .A0(n2348), .A1(n5707), .B0(n2349), .B1(n5678), .C0(n6464), 
        .C1(n5731), .Y(n2351) );
  OAI222XL U8771 ( .A0(n6388), .A1(n5908), .B0(n2311), .B1(n2305), .C0(n367), 
        .C1(n2306), .Y(n4265) );
  AOI211X1 U8772 ( .A0(n5945), .A1(n2307), .B0(n2312), .C0(n5752), .Y(n2311)
         );
  OAI222XL U8773 ( .A0(n2309), .A1(n5707), .B0(n2310), .B1(n5678), .C0(n6465), 
        .C1(n5731), .Y(n2312) );
  OAI222XL U8774 ( .A0(n6389), .A1(n5908), .B0(n2272), .B1(n2266), .C0(n359), 
        .C1(n2267), .Y(n4257) );
  AOI211X1 U8775 ( .A0(n5945), .A1(n2268), .B0(n2273), .C0(n5752), .Y(n2272)
         );
  OAI222XL U8776 ( .A0(n2270), .A1(n5707), .B0(n2271), .B1(n5678), .C0(n6466), 
        .C1(n5731), .Y(n2273) );
  OAI222XL U8777 ( .A0(n6390), .A1(n5908), .B0(n2233), .B1(n2227), .C0(n351), 
        .C1(n2228), .Y(n4249) );
  AOI211X1 U8778 ( .A0(n5945), .A1(n2229), .B0(n2234), .C0(n5752), .Y(n2233)
         );
  OAI222XL U8779 ( .A0(n2231), .A1(n5707), .B0(n2232), .B1(n5678), .C0(n6467), 
        .C1(n5731), .Y(n2234) );
  OAI222XL U8780 ( .A0(n6391), .A1(n5908), .B0(n2194), .B1(n2188), .C0(n343), 
        .C1(n2189), .Y(n4241) );
  AOI211X1 U8781 ( .A0(n5945), .A1(n2190), .B0(n2195), .C0(n5752), .Y(n2194)
         );
  OAI222XL U8782 ( .A0(n2192), .A1(n5707), .B0(n2193), .B1(n5678), .C0(n6468), 
        .C1(n5731), .Y(n2195) );
  OAI222XL U8783 ( .A0(n6392), .A1(n5908), .B0(n2155), .B1(n2149), .C0(n335), 
        .C1(n2150), .Y(n4233) );
  AOI211X1 U8784 ( .A0(n5945), .A1(n2151), .B0(n2156), .C0(n5752), .Y(n2155)
         );
  OAI222XL U8785 ( .A0(n2153), .A1(n5707), .B0(n2154), .B1(n5678), .C0(n6469), 
        .C1(n5731), .Y(n2156) );
  OAI222XL U8786 ( .A0(n6393), .A1(n5908), .B0(n2111), .B1(n2105), .C0(n327), 
        .C1(n2106), .Y(n4225) );
  AOI211X1 U8787 ( .A0(n5945), .A1(n2107), .B0(n2112), .C0(n5752), .Y(n2111)
         );
  OAI222XL U8788 ( .A0(n2109), .A1(n5707), .B0(n2110), .B1(n5678), .C0(n6470), 
        .C1(n5731), .Y(n2112) );
  OAI222XL U8789 ( .A0(n6394), .A1(n5906), .B0(n2072), .B1(n2066), .C0(n319), 
        .C1(n2067), .Y(n4217) );
  AOI211X1 U8790 ( .A0(n5945), .A1(n2068), .B0(n2073), .C0(n5752), .Y(n2072)
         );
  OAI222XL U8791 ( .A0(n2070), .A1(n5706), .B0(n2071), .B1(n5678), .C0(n6471), 
        .C1(n5731), .Y(n2073) );
  OAI222XL U8792 ( .A0(n6395), .A1(n5906), .B0(n2033), .B1(n2027), .C0(n311), 
        .C1(n2028), .Y(n4209) );
  AOI211X1 U8793 ( .A0(n5944), .A1(n2029), .B0(n2034), .C0(n5752), .Y(n2033)
         );
  OAI222XL U8794 ( .A0(n2031), .A1(n5705), .B0(n2032), .B1(n5679), .C0(n6472), 
        .C1(n5731), .Y(n2034) );
  OAI222XL U8795 ( .A0(n6396), .A1(n5906), .B0(n1992), .B1(n1987), .C0(n303), 
        .C1(n1988), .Y(n4201) );
  AOI211X1 U8796 ( .A0(n5944), .A1(n6473), .B0(n1993), .C0(n5752), .Y(n1992)
         );
  OAI222XL U8797 ( .A0(n1990), .A1(n5707), .B0(n1991), .B1(n5679), .C0(n6474), 
        .C1(n5730), .Y(n1993) );
  OAI222XL U8798 ( .A0(n6397), .A1(n5908), .B0(n1953), .B1(n1948), .C0(n295), 
        .C1(n1949), .Y(n4193) );
  AOI211X1 U8799 ( .A0(n5945), .A1(n6475), .B0(n1954), .C0(n5755), .Y(n1953)
         );
  OAI222XL U8800 ( .A0(n1951), .A1(n5706), .B0(n1952), .B1(n5679), .C0(n6476), 
        .C1(n5730), .Y(n1954) );
  OAI222XL U8801 ( .A0(n6398), .A1(n5908), .B0(n1914), .B1(n1909), .C0(n287), 
        .C1(n1910), .Y(n4185) );
  AOI211X1 U8802 ( .A0(n5945), .A1(n6477), .B0(n1915), .C0(n5753), .Y(n1914)
         );
  OAI222XL U8803 ( .A0(n1912), .A1(n5706), .B0(n1913), .B1(n5679), .C0(n6478), 
        .C1(n5730), .Y(n1915) );
  OAI222XL U8804 ( .A0(n4832), .A1(n5907), .B0(n1875), .B1(n1870), .C0(n279), 
        .C1(n1871), .Y(n4177) );
  AOI211X1 U8805 ( .A0(n5944), .A1(n6479), .B0(n1876), .C0(n5754), .Y(n1875)
         );
  OAI222XL U8806 ( .A0(n1873), .A1(n5706), .B0(n1874), .B1(n5679), .C0(n6480), 
        .C1(n5730), .Y(n1876) );
  OAI222XL U8807 ( .A0(n6399), .A1(n5907), .B0(n1836), .B1(n1831), .C0(n271), 
        .C1(n4643), .Y(n4169) );
  AOI211X1 U8808 ( .A0(n5944), .A1(n6481), .B0(n1837), .C0(n5755), .Y(n1836)
         );
  OAI222XL U8809 ( .A0(n1834), .A1(n5707), .B0(n1835), .B1(n5679), .C0(n6482), 
        .C1(n5730), .Y(n1837) );
  OAI222XL U8810 ( .A0(n6400), .A1(n5907), .B0(n1792), .B1(n1787), .C0(n263), 
        .C1(n1788), .Y(n4161) );
  AOI211X1 U8811 ( .A0(n5945), .A1(n6483), .B0(n1793), .C0(n5752), .Y(n1792)
         );
  OAI222XL U8812 ( .A0(n1790), .A1(n5707), .B0(n1791), .B1(n5679), .C0(n6484), 
        .C1(n5730), .Y(n1793) );
  OAI222XL U8813 ( .A0(n6401), .A1(n5906), .B0(n1747), .B1(n1742), .C0(n255), 
        .C1(n1743), .Y(n4153) );
  AOI211X1 U8814 ( .A0(n5944), .A1(n6485), .B0(n1748), .C0(n5753), .Y(n1747)
         );
  OAI222XL U8815 ( .A0(n1745), .A1(n5707), .B0(n1746), .B1(n5679), .C0(n6486), 
        .C1(n5730), .Y(n1748) );
  OAI222XL U8816 ( .A0(n6402), .A1(n5908), .B0(n1703), .B1(n1698), .C0(n247), 
        .C1(n1699), .Y(n4145) );
  AOI211X1 U8817 ( .A0(n5944), .A1(n6487), .B0(n1704), .C0(n5754), .Y(n1703)
         );
  OAI222XL U8818 ( .A0(n1701), .A1(n5706), .B0(n1702), .B1(n5679), .C0(n6488), 
        .C1(n5730), .Y(n1704) );
  OAI222XL U8819 ( .A0(n6403), .A1(n5907), .B0(n1659), .B1(n1654), .C0(n239), 
        .C1(n1655), .Y(n4137) );
  AOI211X1 U8820 ( .A0(n5944), .A1(n6489), .B0(n1660), .C0(n5754), .Y(n1659)
         );
  OAI222XL U8821 ( .A0(n1657), .A1(n5706), .B0(n1658), .B1(n5679), .C0(n6490), 
        .C1(n5730), .Y(n1660) );
  OAI222XL U8822 ( .A0(n6404), .A1(n5907), .B0(n1615), .B1(n1610), .C0(n231), 
        .C1(n1611), .Y(n4129) );
  AOI211X1 U8823 ( .A0(n5945), .A1(n6491), .B0(n1616), .C0(n5752), .Y(n1615)
         );
  OAI222XL U8824 ( .A0(n1613), .A1(n5707), .B0(n1614), .B1(n5679), .C0(n6492), 
        .C1(n5730), .Y(n1616) );
  OAI222XL U8825 ( .A0(n6405), .A1(n5908), .B0(n1571), .B1(n1566), .C0(n223), 
        .C1(n1567), .Y(n4121) );
  AOI211X1 U8826 ( .A0(n5944), .A1(n6493), .B0(n1572), .C0(n5753), .Y(n1571)
         );
  OAI222XL U8827 ( .A0(n1569), .A1(n5705), .B0(n1570), .B1(n5679), .C0(n6494), 
        .C1(n5730), .Y(n1572) );
  OAI222XL U8828 ( .A0(n6406), .A1(n5906), .B0(n1527), .B1(n1522), .C0(n215), 
        .C1(n1523), .Y(n4113) );
  AOI211X1 U8829 ( .A0(n5945), .A1(n6495), .B0(n1528), .C0(n5752), .Y(n1527)
         );
  OAI222XL U8830 ( .A0(n1525), .A1(n5706), .B0(n1526), .B1(n5679), .C0(n6496), 
        .C1(n5730), .Y(n1528) );
  OAI222XL U8831 ( .A0(n6407), .A1(n5908), .B0(n1483), .B1(n1478), .C0(n207), 
        .C1(n1479), .Y(n4105) );
  AOI211X1 U8832 ( .A0(n5944), .A1(n6497), .B0(n1484), .C0(n5754), .Y(n1483)
         );
  OAI222XL U8833 ( .A0(n1481), .A1(n5706), .B0(n1482), .B1(n5680), .C0(n6498), 
        .C1(n5732), .Y(n1484) );
  OAI222XL U8834 ( .A0(n3987), .A1(n5724), .B0(n3988), .B1(n5699), .C0(n6423), 
        .C1(n5750), .Y(n4028) );
  OAI222XL U8835 ( .A0(n3968), .A1(n5863), .B0(n4021), .B1(n3970), .C0(n708), 
        .C1(n6346), .Y(n4606) );
  AOI211X1 U8836 ( .A0(n5921), .A1(n3971), .B0(n4022), .C0(n5861), .Y(n4021)
         );
  OAI222XL U8837 ( .A0(n3987), .A1(n5722), .B0(n3988), .B1(n5695), .C0(n6423), 
        .C1(n5746), .Y(n4022) );
  OAI222XL U8838 ( .A0(n3968), .A1(n5872), .B0(n4015), .B1(n3970), .C0(n707), 
        .C1(n6346), .Y(n4605) );
  OAI222XL U8839 ( .A0(n3987), .A1(n5718), .B0(n3988), .B1(n5691), .C0(n6423), 
        .C1(n5743), .Y(n4016) );
  OAI222XL U8840 ( .A0(n3968), .A1(n5883), .B0(n4009), .B1(n3970), .C0(n706), 
        .C1(n6346), .Y(n4604) );
  AOI211X1 U8841 ( .A0(n5929), .A1(n3971), .B0(n4010), .C0(n5876), .Y(n4009)
         );
  OAI222XL U8842 ( .A0(n3987), .A1(n5716), .B0(n3988), .B1(n5688), .C0(n6423), 
        .C1(n5740), .Y(n4010) );
  AOI211X1 U8843 ( .A0(n5935), .A1(n3971), .B0(n4004), .C0(n5889), .Y(n4003)
         );
  OAI222XL U8844 ( .A0(n3987), .A1(n5711), .B0(n3988), .B1(n5684), .C0(n6423), 
        .C1(n5737), .Y(n4004) );
  OAI222XL U8845 ( .A0(n3968), .A1(n5903), .B0(n3996), .B1(n3970), .C0(n704), 
        .C1(n6346), .Y(n4602) );
  AOI211X1 U8846 ( .A0(n5941), .A1(n3971), .B0(n3997), .C0(n5896), .Y(n3996)
         );
  OAI222XL U8847 ( .A0(n3987), .A1(n6500), .B0(n3988), .B1(n5681), .C0(n6423), 
        .C1(n5735), .Y(n3997) );
  OAI222XL U8848 ( .A0(n3968), .A1(n5909), .B0(n3969), .B1(n3970), .C0(n702), 
        .C1(n6346), .Y(n4600) );
  AOI211X1 U8849 ( .A0(n5948), .A1(n3971), .B0(n3972), .C0(n5759), .Y(n3969)
         );
  OAI222XL U8850 ( .A0(n3987), .A1(n5703), .B0(n3988), .B1(n5675), .C0(n6423), 
        .C1(n5728), .Y(n3972) );
  OAI222XL U8851 ( .A0(n3968), .A1(n5906), .B0(n3989), .B1(n3970), .C0(n703), 
        .C1(n6346), .Y(n4601) );
  AOI211X1 U8852 ( .A0(n5944), .A1(n3971), .B0(n3990), .C0(n5755), .Y(n3989)
         );
  OAI222XL U8853 ( .A0(n3987), .A1(n5705), .B0(n3988), .B1(n5679), .C0(n6423), 
        .C1(n5730), .Y(n3990) );
  MX4X1 U8854 ( .A(n5286), .B(n5284), .C(n5285), .D(n5283), .S0(n5957), .S1(
        n5959), .Y(n5287) );
  MX4X1 U8855 ( .A(\img_buff[24][0] ), .B(\img_buff[25][0] ), .C(
        \img_buff[26][0] ), .D(\img_buff[27][0] ), .S0(n5433), .S1(n5446), .Y(
        n5284) );
  MX4X1 U8856 ( .A(\img_buff[16][0] ), .B(\img_buff[17][0] ), .C(
        \img_buff[18][0] ), .D(\img_buff[19][0] ), .S0(n5434), .S1(n5450), .Y(
        n5286) );
  MX4X1 U8857 ( .A(\img_buff[28][0] ), .B(\img_buff[29][0] ), .C(
        \img_buff[30][0] ), .D(\img_buff[31][0] ), .S0(n5433), .S1(n5446), .Y(
        n5283) );
  MX4X1 U8858 ( .A(n5326), .B(n5324), .C(n5325), .D(n5323), .S0(n4800), .S1(
        n5959), .Y(n5327) );
  MX4X1 U8859 ( .A(\img_buff[16][2] ), .B(\img_buff[17][2] ), .C(
        \img_buff[18][2] ), .D(\img_buff[19][2] ), .S0(n5435), .S1(n4699), .Y(
        n5326) );
  MX4X1 U8860 ( .A(\img_buff[24][2] ), .B(\img_buff[25][2] ), .C(
        \img_buff[26][2] ), .D(\img_buff[27][2] ), .S0(n5435), .S1(n4699), .Y(
        n5324) );
  MX4X1 U8861 ( .A(\img_buff[4][0] ), .B(\img_buff[5][0] ), .C(
        \img_buff[6][0] ), .D(\img_buff[7][0] ), .S0(n5434), .S1(n5450), .Y(
        n5290) );
  MX4X1 U8862 ( .A(\img_buff[52][2] ), .B(\img_buff[53][2] ), .C(
        \img_buff[54][2] ), .D(\img_buff[55][2] ), .S0(n5074), .S1(n5448), .Y(
        n5315) );
  MX4X1 U8863 ( .A(\img_buff[16][3] ), .B(\img_buff[17][3] ), .C(
        \img_buff[18][3] ), .D(\img_buff[19][3] ), .S0(n5436), .S1(n5450), .Y(
        n5346) );
  MX4X1 U8864 ( .A(\img_buff[24][3] ), .B(\img_buff[25][3] ), .C(
        \img_buff[26][3] ), .D(\img_buff[27][3] ), .S0(n5436), .S1(n5450), .Y(
        n5344) );
  MX4X1 U8865 ( .A(\img_buff[28][3] ), .B(\img_buff[29][3] ), .C(
        \img_buff[30][3] ), .D(\img_buff[31][3] ), .S0(n5436), .S1(n5450), .Y(
        n5343) );
  MX4X1 U8866 ( .A(n5366), .B(n5364), .C(n5365), .D(n5363), .S0(n4800), .S1(
        n5959), .Y(n5367) );
  MX4X1 U8867 ( .A(\img_buff[16][4] ), .B(\img_buff[17][4] ), .C(
        \img_buff[18][4] ), .D(\img_buff[19][4] ), .S0(n5436), .S1(n4699), .Y(
        n5366) );
  MX4X1 U8868 ( .A(\img_buff[24][4] ), .B(\img_buff[25][4] ), .C(
        \img_buff[26][4] ), .D(\img_buff[27][4] ), .S0(n5437), .S1(n4699), .Y(
        n5364) );
  MX4X1 U8869 ( .A(\img_buff[28][4] ), .B(\img_buff[29][4] ), .C(
        \img_buff[30][4] ), .D(\img_buff[31][4] ), .S0(n5074), .S1(n4699), .Y(
        n5363) );
  MX4X1 U8870 ( .A(\img_buff[16][5] ), .B(\img_buff[17][5] ), .C(
        \img_buff[18][5] ), .D(\img_buff[19][5] ), .S0(n5438), .S1(n5452), .Y(
        n5386) );
  MX4X1 U8871 ( .A(\img_buff[24][5] ), .B(\img_buff[25][5] ), .C(
        \img_buff[26][5] ), .D(\img_buff[27][5] ), .S0(n5438), .S1(n5452), .Y(
        n5384) );
  MX4X1 U8872 ( .A(\img_buff[16][6] ), .B(\img_buff[17][6] ), .C(
        \img_buff[18][6] ), .D(\img_buff[19][6] ), .S0(n5439), .S1(n5453), .Y(
        n5406) );
  MX4X1 U8873 ( .A(\img_buff[24][6] ), .B(\img_buff[25][6] ), .C(
        \img_buff[26][6] ), .D(\img_buff[27][6] ), .S0(n5439), .S1(n5453), .Y(
        n5404) );
  MX4X1 U8874 ( .A(\img_buff[28][6] ), .B(\img_buff[29][6] ), .C(
        \img_buff[30][6] ), .D(\img_buff[31][6] ), .S0(n5439), .S1(n5453), .Y(
        n5403) );
  MX4X1 U8875 ( .A(\img_buff[20][0] ), .B(\img_buff[21][0] ), .C(
        \img_buff[22][0] ), .D(\img_buff[23][0] ), .S0(n5433), .S1(n5446), .Y(
        n5285) );
  MX4X1 U8876 ( .A(\img_buff[52][0] ), .B(\img_buff[53][0] ), .C(
        \img_buff[54][0] ), .D(\img_buff[55][0] ), .S0(n5433), .S1(n5446), .Y(
        n5275) );
  MX4X1 U8877 ( .A(\img_buff[36][0] ), .B(\img_buff[37][0] ), .C(
        \img_buff[38][0] ), .D(\img_buff[39][0] ), .S0(n5433), .S1(n5446), .Y(
        n5280) );
  MX4X1 U8878 ( .A(\img_buff[0][0] ), .B(\img_buff[1][0] ), .C(
        \img_buff[2][0] ), .D(\img_buff[3][0] ), .S0(n5434), .S1(n5450), .Y(
        n5291) );
  MX4X1 U8879 ( .A(\img_buff[32][2] ), .B(\img_buff[33][2] ), .C(
        \img_buff[34][2] ), .D(\img_buff[35][2] ), .S0(n5435), .S1(n4699), .Y(
        n5321) );
  MX4X1 U8880 ( .A(\img_buff[0][2] ), .B(\img_buff[1][2] ), .C(
        \img_buff[2][2] ), .D(\img_buff[3][2] ), .S0(n5435), .S1(n4699), .Y(
        n5331) );
  MX4X1 U8881 ( .A(\img_buff[32][0] ), .B(\img_buff[33][0] ), .C(
        \img_buff[34][0] ), .D(\img_buff[35][0] ), .S0(n5433), .S1(n5446), .Y(
        n5281) );
  MX4X1 U8882 ( .A(n5276), .B(n5274), .C(n5275), .D(n5273), .S0(n4800), .S1(
        n5959), .Y(n5277) );
  MX4X1 U8883 ( .A(\img_buff[48][0] ), .B(\img_buff[49][0] ), .C(
        \img_buff[50][0] ), .D(\img_buff[51][0] ), .S0(n5433), .S1(n5446), .Y(
        n5276) );
  MX4X1 U8884 ( .A(\img_buff[56][0] ), .B(\img_buff[57][0] ), .C(
        \img_buff[58][0] ), .D(\img_buff[59][0] ), .S0(n5433), .S1(n5446), .Y(
        n5274) );
  MX4X1 U8885 ( .A(\img_buff[60][0] ), .B(\img_buff[61][0] ), .C(
        \img_buff[62][0] ), .D(\img_buff[63][0] ), .S0(n5433), .S1(n5446), .Y(
        n5273) );
  MX4X1 U8886 ( .A(n5316), .B(n5314), .C(n5315), .D(n5313), .S0(n4800), .S1(
        n5959), .Y(n5317) );
  MX4X1 U8887 ( .A(\img_buff[48][2] ), .B(\img_buff[49][2] ), .C(
        \img_buff[50][2] ), .D(\img_buff[51][2] ), .S0(n5433), .S1(n5448), .Y(
        n5316) );
  MX4X1 U8888 ( .A(\img_buff[56][2] ), .B(\img_buff[57][2] ), .C(
        \img_buff[58][2] ), .D(\img_buff[59][2] ), .S0(n5074), .S1(n5448), .Y(
        n5314) );
  MX4X1 U8889 ( .A(\img_buff[60][2] ), .B(\img_buff[61][2] ), .C(
        \img_buff[62][2] ), .D(\img_buff[63][2] ), .S0(n5078), .S1(n5448), .Y(
        n5313) );
  MX4X1 U8890 ( .A(\img_buff[12][0] ), .B(\img_buff[13][0] ), .C(
        \img_buff[14][0] ), .D(\img_buff[15][0] ), .S0(n5434), .S1(n5450), .Y(
        n5288) );
  MX4X1 U8891 ( .A(\img_buff[44][2] ), .B(\img_buff[45][2] ), .C(
        \img_buff[46][2] ), .D(\img_buff[47][2] ), .S0(n5074), .S1(n5448), .Y(
        n5318) );
  MX4X1 U8892 ( .A(\img_buff[48][3] ), .B(\img_buff[49][3] ), .C(
        \img_buff[50][3] ), .D(\img_buff[51][3] ), .S0(n5436), .S1(n5450), .Y(
        n5336) );
  MX4X1 U8893 ( .A(\img_buff[56][3] ), .B(\img_buff[57][3] ), .C(
        \img_buff[58][3] ), .D(\img_buff[59][3] ), .S0(n5435), .S1(n4699), .Y(
        n5334) );
  MX4X1 U8894 ( .A(n5356), .B(n5354), .C(n5355), .D(n5353), .S0(n5957), .S1(
        n5959), .Y(n5357) );
  MX4X1 U8895 ( .A(\img_buff[48][4] ), .B(\img_buff[49][4] ), .C(
        \img_buff[50][4] ), .D(\img_buff[51][4] ), .S0(n5439), .S1(n4699), .Y(
        n5356) );
  MX4X1 U8896 ( .A(\img_buff[56][4] ), .B(\img_buff[57][4] ), .C(
        \img_buff[58][4] ), .D(\img_buff[59][4] ), .S0(n5437), .S1(n5453), .Y(
        n5354) );
  MX4X1 U8897 ( .A(\img_buff[60][4] ), .B(\img_buff[61][4] ), .C(
        \img_buff[62][4] ), .D(\img_buff[63][4] ), .S0(n5436), .S1(n4699), .Y(
        n5353) );
  MX4X1 U8898 ( .A(\img_buff[48][6] ), .B(\img_buff[49][6] ), .C(
        \img_buff[50][6] ), .D(\img_buff[51][6] ), .S0(n5438), .S1(n5452), .Y(
        n5396) );
  MX4X1 U8899 ( .A(\img_buff[56][6] ), .B(\img_buff[57][6] ), .C(
        \img_buff[58][6] ), .D(\img_buff[59][6] ), .S0(n5438), .S1(n5452), .Y(
        n5394) );
  MX4X1 U8900 ( .A(\img_buff[60][6] ), .B(\img_buff[61][6] ), .C(
        \img_buff[62][6] ), .D(\img_buff[63][6] ), .S0(n5438), .S1(n5452), .Y(
        n5393) );
  MX4X1 U8901 ( .A(\img_buff[44][0] ), .B(\img_buff[45][0] ), .C(
        \img_buff[46][0] ), .D(\img_buff[47][0] ), .S0(n5433), .S1(n5446), .Y(
        n5278) );
  MX4X1 U8902 ( .A(\img_buff[8][0] ), .B(\img_buff[9][0] ), .C(
        \img_buff[10][0] ), .D(\img_buff[11][0] ), .S0(n5434), .S1(n5450), .Y(
        n5289) );
  MX4X1 U8903 ( .A(\img_buff[40][2] ), .B(\img_buff[41][2] ), .C(
        \img_buff[42][2] ), .D(\img_buff[43][2] ), .S0(n5435), .S1(n4699), .Y(
        n5319) );
  MX4X1 U8904 ( .A(\img_buff[8][2] ), .B(\img_buff[9][2] ), .C(
        \img_buff[10][2] ), .D(\img_buff[11][2] ), .S0(n5435), .S1(n4699), .Y(
        n5329) );
  MX4X1 U8905 ( .A(\img_buff[40][0] ), .B(\img_buff[41][0] ), .C(
        \img_buff[42][0] ), .D(\img_buff[43][0] ), .S0(n5433), .S1(n5446), .Y(
        n5279) );
  CLKINVX1 U8906 ( .A(n1018), .Y(n6414) );
  AOI222XL U8907 ( .A0(\img_buff[0][0] ), .A1(n6415), .B0(n978), .B1(n1019), 
        .C0(n4884), .C1(n980), .Y(n1018) );
  OAI211X1 U8908 ( .A0(n982), .A1(n5919), .B0(n5796), .C0(n1021), .Y(n1019) );
  AOI222XL U8909 ( .A0(n5666), .A1(n984), .B0(N3351), .B1(n985), .C0(N3359), 
        .C1(n986), .Y(n1021) );
  CLKINVX1 U8910 ( .A(n1013), .Y(n6413) );
  AOI222XL U8911 ( .A0(\img_buff[0][1] ), .A1(n6415), .B0(n978), .B1(n1014), 
        .C0(n4885), .C1(n980), .Y(n1013) );
  OAI211X1 U8912 ( .A0(n982), .A1(n5924), .B0(n5862), .C0(n1016), .Y(n1014) );
  AOI222XL U8913 ( .A0(n5665), .A1(n984), .B0(n5657), .B1(n985), .C0(N3358), 
        .C1(n986), .Y(n1016) );
  CLKINVX1 U8914 ( .A(n1008), .Y(n6412) );
  AOI222XL U8915 ( .A0(\img_buff[0][2] ), .A1(n6415), .B0(n978), .B1(n1009), 
        .C0(n4886), .C1(n980), .Y(n1008) );
  OAI211X1 U8916 ( .A0(n982), .A1(n5927), .B0(n5870), .C0(n1011), .Y(n1009) );
  AOI222XL U8917 ( .A0(n5664), .A1(n984), .B0(n5656), .B1(n985), .C0(N3357), 
        .C1(n986), .Y(n1011) );
  CLKINVX1 U8918 ( .A(n1003), .Y(n6411) );
  AOI222XL U8919 ( .A0(\img_buff[0][3] ), .A1(n6415), .B0(n978), .B1(n1004), 
        .C0(n4887), .C1(n980), .Y(n1003) );
  OAI211X1 U8920 ( .A0(n982), .A1(n5931), .B0(n5882), .C0(n1006), .Y(n1004) );
  AOI222XL U8921 ( .A0(n5663), .A1(n984), .B0(n5655), .B1(n985), .C0(n4667), 
        .C1(n986), .Y(n1006) );
  CLKINVX1 U8922 ( .A(n998), .Y(n6410) );
  AOI222XL U8923 ( .A0(\img_buff[0][4] ), .A1(n6415), .B0(n978), .B1(n999), 
        .C0(n4888), .C1(n980), .Y(n998) );
  OAI211X1 U8924 ( .A0(n982), .A1(n5938), .B0(n5890), .C0(n1001), .Y(n999) );
  AOI222XL U8925 ( .A0(n5662), .A1(n984), .B0(n5654), .B1(n985), .C0(N3355), 
        .C1(n986), .Y(n1001) );
  CLKINVX1 U8926 ( .A(n993), .Y(n6409) );
  AOI222XL U8927 ( .A0(\img_buff[0][5] ), .A1(n6415), .B0(n978), .B1(n994), 
        .C0(n4889), .C1(n980), .Y(n993) );
  OAI211X1 U8928 ( .A0(n982), .A1(n5943), .B0(n5902), .C0(n996), .Y(n994) );
  AOI222XL U8929 ( .A0(n5661), .A1(n984), .B0(n5653), .B1(n985), .C0(n5659), 
        .C1(n986), .Y(n996) );
  CLKINVX1 U8930 ( .A(n977), .Y(n6408) );
  AOI222XL U8931 ( .A0(\img_buff[0][7] ), .A1(n6415), .B0(n978), .B1(n979), 
        .C0(n4890), .C1(n980), .Y(n977) );
  OAI211X1 U8932 ( .A0(n982), .A1(n5950), .B0(n4669), .C0(n983), .Y(n979) );
  AOI222XL U8933 ( .A0(N3360), .A1(n984), .B0(n5651), .B1(n985), .C0(n5658), 
        .C1(n986), .Y(n983) );
  OAI211XL U8934 ( .A0(n982), .A1(n5946), .B0(n4814), .C0(n991), .Y(n989) );
  AOI222XL U8935 ( .A0(n5660), .A1(n984), .B0(n5652), .B1(n985), .C0(N3353), 
        .C1(n986), .Y(n991) );
  MX4X1 U8936 ( .A(\img_buff[24][0] ), .B(\img_buff[25][0] ), .C(
        \img_buff[26][0] ), .D(\img_buff[27][0] ), .S0(n5245), .S1(n5639), .Y(
        n5475) );
  MX4X1 U8937 ( .A(\img_buff[28][0] ), .B(\img_buff[29][0] ), .C(
        \img_buff[30][0] ), .D(\img_buff[31][0] ), .S0(n5244), .S1(n5639), .Y(
        n5474) );
  MX4X1 U8938 ( .A(\img_buff[20][0] ), .B(\img_buff[21][0] ), .C(
        \img_buff[22][0] ), .D(\img_buff[23][0] ), .S0(n5624), .S1(n5639), .Y(
        n5476) );
  MX4X1 U8939 ( .A(n5497), .B(n5495), .C(n5496), .D(n5494), .S0(n5648), .S1(
        n5269), .Y(n5498) );
  MX4X1 U8940 ( .A(\img_buff[4][0] ), .B(\img_buff[5][0] ), .C(
        \img_buff[6][0] ), .D(\img_buff[7][0] ), .S0(n5628), .S1(n5640), .Y(
        n5481) );
  MX4X1 U8941 ( .A(\img_buff[20][2] ), .B(\img_buff[21][2] ), .C(
        \img_buff[22][2] ), .D(\img_buff[23][2] ), .S0(n5629), .S1(n5266), .Y(
        n5516) );
  MX4X1 U8942 ( .A(\img_buff[52][2] ), .B(\img_buff[53][2] ), .C(
        \img_buff[54][2] ), .D(\img_buff[55][2] ), .S0(n5626), .S1(n5641), .Y(
        n5506) );
  MX4X1 U8943 ( .A(\img_buff[36][2] ), .B(\img_buff[37][2] ), .C(
        \img_buff[38][2] ), .D(\img_buff[39][2] ), .S0(n5629), .S1(n5266), .Y(
        n5511) );
  MX4X1 U8944 ( .A(\img_buff[4][2] ), .B(\img_buff[5][2] ), .C(
        \img_buff[6][2] ), .D(\img_buff[7][2] ), .S0(n5629), .S1(n5256), .Y(
        n5521) );
  MX4X1 U8945 ( .A(\img_buff[4][4] ), .B(\img_buff[5][4] ), .C(
        \img_buff[6][4] ), .D(\img_buff[7][4] ), .S0(n5632), .S1(n5644), .Y(
        n5561) );
  MX4X1 U8946 ( .A(\img_buff[4][0] ), .B(\img_buff[5][0] ), .C(
        \img_buff[6][0] ), .D(\img_buff[7][0] ), .S0(n5248), .S1(n5257), .Y(
        n5100) );
  MX4X1 U8947 ( .A(n5517), .B(n5515), .C(n5516), .D(n5514), .S0(n5648), .S1(
        n5269), .Y(n5518) );
  MX4X1 U8948 ( .A(\img_buff[16][2] ), .B(\img_buff[17][2] ), .C(
        \img_buff[18][2] ), .D(\img_buff[19][2] ), .S0(n5629), .S1(n4749), .Y(
        n5517) );
  MX4X1 U8949 ( .A(\img_buff[24][2] ), .B(\img_buff[25][2] ), .C(
        \img_buff[26][2] ), .D(\img_buff[27][2] ), .S0(n5629), .S1(n5259), .Y(
        n5515) );
  MX4X1 U8950 ( .A(\img_buff[28][2] ), .B(\img_buff[29][2] ), .C(
        \img_buff[30][2] ), .D(\img_buff[31][2] ), .S0(n5629), .S1(n5256), .Y(
        n5514) );
  MX4X1 U8951 ( .A(\img_buff[20][2] ), .B(\img_buff[21][2] ), .C(
        \img_buff[22][2] ), .D(\img_buff[23][2] ), .S0(n5250), .S1(n5259), .Y(
        n5135) );
  MX4X1 U8952 ( .A(\img_buff[52][2] ), .B(\img_buff[53][2] ), .C(
        \img_buff[54][2] ), .D(\img_buff[55][2] ), .S0(n5249), .S1(n5258), .Y(
        n5125) );
  MX4X1 U8953 ( .A(\img_buff[36][2] ), .B(\img_buff[37][2] ), .C(
        \img_buff[38][2] ), .D(\img_buff[39][2] ), .S0(n5250), .S1(n5259), .Y(
        n5130) );
  MX4X1 U8954 ( .A(\img_buff[4][2] ), .B(\img_buff[5][2] ), .C(
        \img_buff[6][2] ), .D(\img_buff[7][2] ), .S0(n5250), .S1(n5259), .Y(
        n5140) );
  MX4X1 U8955 ( .A(\img_buff[20][3] ), .B(\img_buff[21][3] ), .C(
        \img_buff[22][3] ), .D(\img_buff[23][3] ), .S0(n5436), .S1(n5450), .Y(
        n5345) );
  MX4X1 U8956 ( .A(\img_buff[52][3] ), .B(\img_buff[53][3] ), .C(
        \img_buff[54][3] ), .D(\img_buff[55][3] ), .S0(n5436), .S1(n5450), .Y(
        n5335) );
  MX4X1 U8957 ( .A(\img_buff[36][3] ), .B(\img_buff[37][3] ), .C(
        \img_buff[38][3] ), .D(\img_buff[39][3] ), .S0(n5436), .S1(n5450), .Y(
        n5340) );
  MX4X1 U8958 ( .A(\img_buff[4][3] ), .B(\img_buff[5][3] ), .C(
        \img_buff[6][3] ), .D(\img_buff[7][3] ), .S0(n5436), .S1(n5450), .Y(
        n5350) );
  MX4X1 U8959 ( .A(\img_buff[20][4] ), .B(\img_buff[21][4] ), .C(
        \img_buff[22][4] ), .D(\img_buff[23][4] ), .S0(n5434), .S1(n5453), .Y(
        n5365) );
  MX4X1 U8960 ( .A(\img_buff[52][4] ), .B(\img_buff[53][4] ), .C(
        \img_buff[54][4] ), .D(\img_buff[55][4] ), .S0(n5076), .S1(n5453), .Y(
        n5355) );
  MX4X1 U8961 ( .A(\img_buff[36][4] ), .B(\img_buff[37][4] ), .C(
        \img_buff[38][4] ), .D(\img_buff[39][4] ), .S0(n5433), .S1(n4699), .Y(
        n5360) );
  MX4X1 U8962 ( .A(\img_buff[4][4] ), .B(\img_buff[5][4] ), .C(
        \img_buff[6][4] ), .D(\img_buff[7][4] ), .S0(n5437), .S1(n5451), .Y(
        n5370) );
  MX4X1 U8963 ( .A(\img_buff[20][4] ), .B(\img_buff[21][4] ), .C(
        \img_buff[22][4] ), .D(\img_buff[23][4] ), .S0(n5077), .S1(n5058), .Y(
        n4987) );
  MX4X1 U8964 ( .A(\img_buff[52][4] ), .B(\img_buff[53][4] ), .C(
        \img_buff[54][4] ), .D(\img_buff[55][4] ), .S0(n5077), .S1(n5064), .Y(
        n4977) );
  MX4X1 U8965 ( .A(\img_buff[36][4] ), .B(\img_buff[37][4] ), .C(
        \img_buff[38][4] ), .D(\img_buff[39][4] ), .S0(n5077), .S1(n5055), .Y(
        n4982) );
  MX4X1 U8966 ( .A(\img_buff[4][4] ), .B(\img_buff[5][4] ), .C(
        \img_buff[6][4] ), .D(\img_buff[7][4] ), .S0(n5078), .S1(n5056), .Y(
        n4992) );
  MX4X1 U8967 ( .A(\img_buff[20][5] ), .B(\img_buff[21][5] ), .C(
        \img_buff[22][5] ), .D(\img_buff[23][5] ), .S0(n5438), .S1(n5452), .Y(
        n5385) );
  MX4X1 U8968 ( .A(\img_buff[4][5] ), .B(\img_buff[5][5] ), .C(
        \img_buff[6][5] ), .D(\img_buff[7][5] ), .S0(n5438), .S1(n5452), .Y(
        n5390) );
  MX4X1 U8969 ( .A(\img_buff[20][6] ), .B(\img_buff[21][6] ), .C(
        \img_buff[22][6] ), .D(\img_buff[23][6] ), .S0(n5439), .S1(n5453), .Y(
        n5405) );
  MX4X1 U8970 ( .A(\img_buff[52][6] ), .B(\img_buff[53][6] ), .C(
        \img_buff[54][6] ), .D(\img_buff[55][6] ), .S0(n5438), .S1(n5452), .Y(
        n5395) );
  MX4X1 U8971 ( .A(\img_buff[36][6] ), .B(\img_buff[37][6] ), .C(
        \img_buff[38][6] ), .D(\img_buff[39][6] ), .S0(n5439), .S1(n5453), .Y(
        n5400) );
  MX4X1 U8972 ( .A(\img_buff[4][6] ), .B(\img_buff[5][6] ), .C(
        \img_buff[6][6] ), .D(\img_buff[7][6] ), .S0(n5439), .S1(n5453), .Y(
        n5410) );
  MX4X1 U8973 ( .A(n5096), .B(n5094), .C(n5095), .D(n5093), .S0(n5272), .S1(
        n5647), .Y(n5097) );
  MX4X1 U8974 ( .A(\img_buff[24][0] ), .B(\img_buff[25][0] ), .C(
        \img_buff[26][0] ), .D(\img_buff[27][0] ), .S0(n4653), .S1(n5644), .Y(
        n5094) );
  MX4X1 U8975 ( .A(\img_buff[28][0] ), .B(\img_buff[29][0] ), .C(
        \img_buff[30][0] ), .D(\img_buff[31][0] ), .S0(n4653), .S1(n5266), .Y(
        n5093) );
  MX4X1 U8976 ( .A(\img_buff[20][0] ), .B(\img_buff[21][0] ), .C(
        \img_buff[22][0] ), .D(\img_buff[23][0] ), .S0(n4653), .S1(n5641), .Y(
        n5095) );
  MX4X1 U8977 ( .A(n4928), .B(n4926), .C(n4927), .D(n4925), .S0(n5068), .S1(
        n5969), .Y(n4929) );
  MX4X1 U8978 ( .A(\img_buff[28][1] ), .B(\img_buff[29][1] ), .C(
        \img_buff[30][1] ), .D(\img_buff[31][1] ), .S0(n5436), .S1(n5058), .Y(
        n4925) );
  MX4X1 U8979 ( .A(\img_buff[20][1] ), .B(\img_buff[21][1] ), .C(
        \img_buff[22][1] ), .D(\img_buff[23][1] ), .S0(n5436), .S1(n4762), .Y(
        n4927) );
  MX4X1 U8980 ( .A(\img_buff[24][1] ), .B(\img_buff[25][1] ), .C(
        \img_buff[26][1] ), .D(\img_buff[27][1] ), .S0(n5436), .S1(n5057), .Y(
        n4926) );
  MX4X1 U8981 ( .A(n5136), .B(n5134), .C(n5135), .D(n5133), .S0(n5272), .S1(
        n5267), .Y(n5137) );
  MX4X1 U8982 ( .A(\img_buff[16][2] ), .B(\img_buff[17][2] ), .C(
        \img_buff[18][2] ), .D(\img_buff[19][2] ), .S0(n5250), .S1(n5259), .Y(
        n5136) );
  MX4X1 U8983 ( .A(\img_buff[24][2] ), .B(\img_buff[25][2] ), .C(
        \img_buff[26][2] ), .D(\img_buff[27][2] ), .S0(n5250), .S1(n5259), .Y(
        n5134) );
  MX4X1 U8984 ( .A(\img_buff[28][2] ), .B(\img_buff[29][2] ), .C(
        \img_buff[30][2] ), .D(\img_buff[31][2] ), .S0(n5250), .S1(n5259), .Y(
        n5133) );
  MX4X1 U8985 ( .A(n4988), .B(n4986), .C(n4987), .D(n4985), .S0(n5068), .S1(
        n5969), .Y(n4989) );
  MX4X1 U8986 ( .A(\img_buff[16][4] ), .B(\img_buff[17][4] ), .C(
        \img_buff[18][4] ), .D(\img_buff[19][4] ), .S0(n5077), .S1(n5061), .Y(
        n4988) );
  MX4X1 U8987 ( .A(\img_buff[24][4] ), .B(\img_buff[25][4] ), .C(
        \img_buff[26][4] ), .D(\img_buff[27][4] ), .S0(n5077), .S1(n5056), .Y(
        n4986) );
  MX4X1 U8988 ( .A(\img_buff[28][4] ), .B(\img_buff[29][4] ), .C(
        \img_buff[30][4] ), .D(\img_buff[31][4] ), .S0(n5077), .S1(n5059), .Y(
        n4985) );
  MX4X1 U8989 ( .A(\img_buff[16][6] ), .B(\img_buff[17][6] ), .C(
        \img_buff[18][6] ), .D(\img_buff[19][6] ), .S0(n5080), .S1(n4762), .Y(
        n5028) );
  MX4X1 U8990 ( .A(\img_buff[24][6] ), .B(\img_buff[25][6] ), .C(
        \img_buff[26][6] ), .D(\img_buff[27][6] ), .S0(n5080), .S1(n5058), .Y(
        n5026) );
  MX4X1 U8991 ( .A(\img_buff[28][6] ), .B(\img_buff[29][6] ), .C(
        \img_buff[30][6] ), .D(\img_buff[31][6] ), .S0(n5080), .S1(n5059), .Y(
        n5025) );
  MX4X1 U8992 ( .A(\img_buff[52][0] ), .B(\img_buff[53][0] ), .C(
        \img_buff[54][0] ), .D(\img_buff[55][0] ), .S0(n5245), .S1(n5639), .Y(
        n5466) );
  MX4X1 U8993 ( .A(\img_buff[36][0] ), .B(\img_buff[37][0] ), .C(
        \img_buff[38][0] ), .D(\img_buff[39][0] ), .S0(n5245), .S1(n5639), .Y(
        n5471) );
  MX4X1 U8994 ( .A(\img_buff[20][0] ), .B(\img_buff[21][0] ), .C(
        \img_buff[22][0] ), .D(\img_buff[23][0] ), .S0(n5073), .S1(n5063), .Y(
        n4907) );
  MX4X1 U8995 ( .A(\img_buff[52][0] ), .B(\img_buff[53][0] ), .C(
        \img_buff[54][0] ), .D(\img_buff[55][0] ), .S0(n5073), .S1(n5056), .Y(
        n4897) );
  MX4X1 U8996 ( .A(\img_buff[52][0] ), .B(\img_buff[53][0] ), .C(
        \img_buff[54][0] ), .D(\img_buff[55][0] ), .S0(n4653), .S1(n5641), .Y(
        n5085) );
  MX4X1 U8997 ( .A(\img_buff[36][0] ), .B(\img_buff[37][0] ), .C(
        \img_buff[38][0] ), .D(\img_buff[39][0] ), .S0(n4653), .S1(n5266), .Y(
        n5090) );
  MX4X1 U8998 ( .A(n5482), .B(n5480), .C(n5481), .D(n5479), .S0(n5649), .S1(
        n5647), .Y(n5483) );
  MX4X1 U8999 ( .A(\img_buff[0][0] ), .B(\img_buff[1][0] ), .C(
        \img_buff[2][0] ), .D(\img_buff[3][0] ), .S0(n5628), .S1(n5640), .Y(
        n5482) );
  MX4X1 U9000 ( .A(\img_buff[8][0] ), .B(\img_buff[9][0] ), .C(
        \img_buff[10][0] ), .D(\img_buff[11][0] ), .S0(n5628), .S1(n5640), .Y(
        n5480) );
  MX4X1 U9001 ( .A(\img_buff[12][0] ), .B(\img_buff[13][0] ), .C(
        \img_buff[14][0] ), .D(\img_buff[15][0] ), .S0(n5628), .S1(n5640), .Y(
        n5479) );
  MX4X1 U9002 ( .A(n4913), .B(n4911), .C(n4912), .D(n4910), .S0(n5067), .S1(
        n5065), .Y(n4914) );
  MX4X1 U9003 ( .A(\img_buff[12][0] ), .B(\img_buff[13][0] ), .C(
        \img_buff[14][0] ), .D(\img_buff[15][0] ), .S0(n5074), .S1(n5060), .Y(
        n4910) );
  MX4X1 U9004 ( .A(\img_buff[4][0] ), .B(\img_buff[5][0] ), .C(
        \img_buff[6][0] ), .D(\img_buff[7][0] ), .S0(n5074), .S1(n5064), .Y(
        n4912) );
  MX4X1 U9005 ( .A(\img_buff[8][0] ), .B(\img_buff[9][0] ), .C(
        \img_buff[10][0] ), .D(\img_buff[11][0] ), .S0(n5074), .S1(n5055), .Y(
        n4911) );
  MX4X1 U9006 ( .A(\img_buff[0][2] ), .B(\img_buff[1][2] ), .C(
        \img_buff[2][2] ), .D(\img_buff[3][2] ), .S0(n5629), .S1(n5256), .Y(
        n5522) );
  MX4X1 U9007 ( .A(\img_buff[0][4] ), .B(\img_buff[1][4] ), .C(
        \img_buff[2][4] ), .D(\img_buff[3][4] ), .S0(n5632), .S1(n5644), .Y(
        n5562) );
  MX4X1 U9008 ( .A(\img_buff[0][0] ), .B(\img_buff[1][0] ), .C(
        \img_buff[2][0] ), .D(\img_buff[3][0] ), .S0(n5074), .S1(n4631), .Y(
        n4913) );
  MX4X1 U9009 ( .A(\img_buff[16][0] ), .B(\img_buff[17][0] ), .C(
        \img_buff[18][0] ), .D(\img_buff[19][0] ), .S0(n5074), .S1(n5970), .Y(
        n4908) );
  MX4X1 U9010 ( .A(\img_buff[16][0] ), .B(\img_buff[17][0] ), .C(
        \img_buff[18][0] ), .D(\img_buff[19][0] ), .S0(n5248), .S1(n5257), .Y(
        n5096) );
  MX4X1 U9011 ( .A(\img_buff[32][2] ), .B(\img_buff[33][2] ), .C(
        \img_buff[34][2] ), .D(\img_buff[35][2] ), .S0(n5250), .S1(n5259), .Y(
        n5131) );
  MX4X1 U9012 ( .A(\img_buff[0][2] ), .B(\img_buff[1][2] ), .C(
        \img_buff[2][2] ), .D(\img_buff[3][2] ), .S0(n5250), .S1(n5259), .Y(
        n5141) );
  MX4X1 U9013 ( .A(\img_buff[32][3] ), .B(\img_buff[33][3] ), .C(
        \img_buff[34][3] ), .D(\img_buff[35][3] ), .S0(n5436), .S1(n5450), .Y(
        n5341) );
  MX4X1 U9014 ( .A(\img_buff[32][4] ), .B(\img_buff[33][4] ), .C(
        \img_buff[34][4] ), .D(\img_buff[35][4] ), .S0(n5435), .S1(n4699), .Y(
        n5361) );
  MX4X1 U9015 ( .A(\img_buff[0][4] ), .B(\img_buff[1][4] ), .C(
        \img_buff[2][4] ), .D(\img_buff[3][4] ), .S0(n5437), .S1(n5451), .Y(
        n5371) );
  MX4X1 U9016 ( .A(\img_buff[32][4] ), .B(\img_buff[33][4] ), .C(
        \img_buff[34][4] ), .D(\img_buff[35][4] ), .S0(n5077), .S1(n4632), .Y(
        n4983) );
  MX4X1 U9017 ( .A(\img_buff[0][4] ), .B(\img_buff[1][4] ), .C(
        \img_buff[2][4] ), .D(\img_buff[3][4] ), .S0(n5078), .S1(n5970), .Y(
        n4993) );
  MX4X1 U9018 ( .A(\img_buff[0][5] ), .B(\img_buff[1][5] ), .C(
        \img_buff[2][5] ), .D(\img_buff[3][5] ), .S0(n5438), .S1(n5452), .Y(
        n5391) );
  MX4X1 U9019 ( .A(\img_buff[32][6] ), .B(\img_buff[33][6] ), .C(
        \img_buff[34][6] ), .D(\img_buff[35][6] ), .S0(n5439), .S1(n5453), .Y(
        n5401) );
  MX4X1 U9020 ( .A(\img_buff[0][6] ), .B(\img_buff[1][6] ), .C(
        \img_buff[2][6] ), .D(\img_buff[3][6] ), .S0(n5439), .S1(n5453), .Y(
        n5411) );
  MX4X1 U9021 ( .A(n5101), .B(n5099), .C(n5100), .D(n5098), .S0(n5272), .S1(
        n5267), .Y(n5102) );
  MX4X1 U9022 ( .A(\img_buff[0][0] ), .B(\img_buff[1][0] ), .C(
        \img_buff[2][0] ), .D(\img_buff[3][0] ), .S0(n5248), .S1(n5257), .Y(
        n5101) );
  MX4X1 U9023 ( .A(\img_buff[8][0] ), .B(\img_buff[9][0] ), .C(
        \img_buff[10][0] ), .D(\img_buff[11][0] ), .S0(n5248), .S1(n5257), .Y(
        n5099) );
  MX4X1 U9024 ( .A(\img_buff[12][0] ), .B(\img_buff[13][0] ), .C(
        \img_buff[14][0] ), .D(\img_buff[15][0] ), .S0(n5248), .S1(n5257), .Y(
        n5098) );
  MX4X1 U9025 ( .A(n4933), .B(n4931), .C(n4932), .D(n4930), .S0(n5068), .S1(
        n5969), .Y(n4934) );
  MX4X1 U9026 ( .A(\img_buff[12][1] ), .B(\img_buff[13][1] ), .C(
        \img_buff[14][1] ), .D(\img_buff[15][1] ), .S0(n5439), .S1(n5061), .Y(
        n4930) );
  MX4X1 U9027 ( .A(\img_buff[4][1] ), .B(\img_buff[5][1] ), .C(
        \img_buff[6][1] ), .D(\img_buff[7][1] ), .S0(n5436), .S1(n5055), .Y(
        n4932) );
  MX4X1 U9028 ( .A(\img_buff[8][1] ), .B(\img_buff[9][1] ), .C(
        \img_buff[10][1] ), .D(\img_buff[11][1] ), .S0(n5436), .S1(n5055), .Y(
        n4931) );
  MX4X1 U9029 ( .A(\img_buff[12][3] ), .B(\img_buff[13][3] ), .C(
        \img_buff[14][3] ), .D(\img_buff[15][3] ), .S0(n5076), .S1(n5060), .Y(
        n4970) );
  MX4X1 U9030 ( .A(\img_buff[4][3] ), .B(\img_buff[5][3] ), .C(
        \img_buff[6][3] ), .D(\img_buff[7][3] ), .S0(n5076), .S1(n5060), .Y(
        n4972) );
  MX4X1 U9031 ( .A(\img_buff[12][7] ), .B(\img_buff[13][7] ), .C(
        \img_buff[14][7] ), .D(\img_buff[15][7] ), .S0(n5440), .S1(n5454), .Y(
        n5428) );
  MX4X1 U9032 ( .A(\img_buff[4][7] ), .B(\img_buff[5][7] ), .C(
        \img_buff[6][7] ), .D(\img_buff[7][7] ), .S0(n5440), .S1(n5454), .Y(
        n5430) );
  MX4X1 U9033 ( .A(\img_buff[8][7] ), .B(\img_buff[9][7] ), .C(
        \img_buff[10][7] ), .D(\img_buff[11][7] ), .S0(n5440), .S1(n5454), .Y(
        n5429) );
  MX4X1 U9034 ( .A(\img_buff[32][0] ), .B(\img_buff[33][0] ), .C(
        \img_buff[34][0] ), .D(\img_buff[35][0] ), .S0(n5254), .S1(n5639), .Y(
        n5472) );
  MX4X1 U9035 ( .A(\img_buff[32][0] ), .B(\img_buff[33][0] ), .C(
        \img_buff[34][0] ), .D(\img_buff[35][0] ), .S0(n5073), .S1(n5064), .Y(
        n4903) );
  MX4X1 U9036 ( .A(\img_buff[48][0] ), .B(\img_buff[49][0] ), .C(
        \img_buff[50][0] ), .D(\img_buff[51][0] ), .S0(n5073), .S1(n5057), .Y(
        n4898) );
  MX4X1 U9037 ( .A(\img_buff[48][0] ), .B(\img_buff[49][0] ), .C(
        \img_buff[50][0] ), .D(\img_buff[51][0] ), .S0(n4653), .S1(n5641), .Y(
        n5086) );
  MX4X1 U9038 ( .A(\img_buff[32][0] ), .B(\img_buff[33][0] ), .C(
        \img_buff[34][0] ), .D(\img_buff[35][0] ), .S0(n4653), .S1(n5641), .Y(
        n5091) );
  MX4X1 U9039 ( .A(n5467), .B(n5465), .C(n5466), .D(n5464), .S0(n5649), .S1(
        n5647), .Y(n5468) );
  MX4X1 U9040 ( .A(\img_buff[48][0] ), .B(\img_buff[49][0] ), .C(
        \img_buff[50][0] ), .D(\img_buff[51][0] ), .S0(n5245), .S1(n5639), .Y(
        n5467) );
  MX4X1 U9041 ( .A(\img_buff[56][0] ), .B(\img_buff[57][0] ), .C(
        \img_buff[58][0] ), .D(\img_buff[59][0] ), .S0(n5243), .S1(n5639), .Y(
        n5465) );
  MX4X1 U9042 ( .A(\img_buff[60][0] ), .B(\img_buff[61][0] ), .C(
        \img_buff[62][0] ), .D(\img_buff[63][0] ), .S0(n5624), .S1(n5639), .Y(
        n5464) );
  MX4X1 U9043 ( .A(\img_buff[12][2] ), .B(\img_buff[13][2] ), .C(
        \img_buff[14][2] ), .D(\img_buff[15][2] ), .S0(n5629), .S1(n5259), .Y(
        n5519) );
  MX4X1 U9044 ( .A(\img_buff[12][4] ), .B(\img_buff[13][4] ), .C(
        \img_buff[14][4] ), .D(\img_buff[15][4] ), .S0(n5632), .S1(n5644), .Y(
        n5559) );
  MX4X1 U9045 ( .A(n5507), .B(n5505), .C(n5506), .D(n5504), .S0(n5648), .S1(
        n5269), .Y(n5508) );
  MX4X1 U9046 ( .A(\img_buff[48][2] ), .B(\img_buff[49][2] ), .C(
        \img_buff[50][2] ), .D(\img_buff[51][2] ), .S0(n5626), .S1(n5641), .Y(
        n5507) );
  MX4X1 U9047 ( .A(\img_buff[56][2] ), .B(\img_buff[57][2] ), .C(
        \img_buff[58][2] ), .D(\img_buff[59][2] ), .S0(n5626), .S1(n5641), .Y(
        n5505) );
  MX4X1 U9048 ( .A(\img_buff[60][2] ), .B(\img_buff[61][2] ), .C(
        \img_buff[62][2] ), .D(\img_buff[63][2] ), .S0(n5626), .S1(n5641), .Y(
        n5504) );
  MX4X1 U9049 ( .A(\img_buff[44][2] ), .B(\img_buff[45][2] ), .C(
        \img_buff[46][2] ), .D(\img_buff[47][2] ), .S0(n5249), .S1(n5258), .Y(
        n5128) );
  MX4X1 U9050 ( .A(\img_buff[12][2] ), .B(\img_buff[13][2] ), .C(
        \img_buff[14][2] ), .D(\img_buff[15][2] ), .S0(n5250), .S1(n5259), .Y(
        n5138) );
  MX4X1 U9051 ( .A(\img_buff[44][3] ), .B(\img_buff[45][3] ), .C(
        \img_buff[46][3] ), .D(\img_buff[47][3] ), .S0(n5436), .S1(n5450), .Y(
        n5338) );
  MX4X1 U9052 ( .A(\img_buff[12][3] ), .B(\img_buff[13][3] ), .C(
        \img_buff[14][3] ), .D(\img_buff[15][3] ), .S0(n5436), .S1(n5450), .Y(
        n5348) );
  MX4X1 U9053 ( .A(n5547), .B(n5545), .C(n5546), .D(n5544), .S0(n5648), .S1(
        n5647), .Y(n5548) );
  MX4X1 U9054 ( .A(\img_buff[44][4] ), .B(\img_buff[45][4] ), .C(
        \img_buff[46][4] ), .D(\img_buff[47][4] ), .S0(n5434), .S1(n4699), .Y(
        n5358) );
  MX4X1 U9055 ( .A(\img_buff[12][4] ), .B(\img_buff[13][4] ), .C(
        \img_buff[14][4] ), .D(\img_buff[15][4] ), .S0(n5437), .S1(n5451), .Y(
        n5368) );
  MX4X1 U9056 ( .A(\img_buff[44][4] ), .B(\img_buff[45][4] ), .C(
        \img_buff[46][4] ), .D(\img_buff[47][4] ), .S0(n5077), .S1(n5059), .Y(
        n4980) );
  MX4X1 U9057 ( .A(\img_buff[12][4] ), .B(\img_buff[13][4] ), .C(
        \img_buff[14][4] ), .D(\img_buff[15][4] ), .S0(n5078), .S1(n5061), .Y(
        n4990) );
  MX4X1 U9058 ( .A(\img_buff[12][5] ), .B(\img_buff[13][5] ), .C(
        \img_buff[14][5] ), .D(\img_buff[15][5] ), .S0(n5438), .S1(n5452), .Y(
        n5388) );
  MX4X1 U9059 ( .A(\img_buff[44][6] ), .B(\img_buff[45][6] ), .C(
        \img_buff[46][6] ), .D(\img_buff[47][6] ), .S0(n5438), .S1(n5452), .Y(
        n5398) );
  MX4X1 U9060 ( .A(\img_buff[12][6] ), .B(\img_buff[13][6] ), .C(
        \img_buff[14][6] ), .D(\img_buff[15][6] ), .S0(n5439), .S1(n5453), .Y(
        n5408) );
  MX4X1 U9061 ( .A(n5126), .B(n5124), .C(n5125), .D(n5123), .S0(n5272), .S1(
        n5267), .Y(n5127) );
  MX4X1 U9062 ( .A(\img_buff[48][2] ), .B(\img_buff[49][2] ), .C(
        \img_buff[50][2] ), .D(\img_buff[51][2] ), .S0(n5249), .S1(n5258), .Y(
        n5126) );
  MX4X1 U9063 ( .A(\img_buff[56][2] ), .B(\img_buff[57][2] ), .C(
        \img_buff[58][2] ), .D(\img_buff[59][2] ), .S0(n5249), .S1(n5258), .Y(
        n5124) );
  MX4X1 U9064 ( .A(\img_buff[60][2] ), .B(\img_buff[61][2] ), .C(
        \img_buff[62][2] ), .D(\img_buff[63][2] ), .S0(n5249), .S1(n5258), .Y(
        n5123) );
  MX4X1 U9065 ( .A(n4978), .B(n4976), .C(n4977), .D(n4975), .S0(n5068), .S1(
        n5969), .Y(n4979) );
  MX4X1 U9066 ( .A(\img_buff[48][4] ), .B(\img_buff[49][4] ), .C(
        \img_buff[50][4] ), .D(\img_buff[51][4] ), .S0(n5077), .S1(n5056), .Y(
        n4978) );
  MX4X1 U9067 ( .A(\img_buff[56][4] ), .B(\img_buff[57][4] ), .C(
        \img_buff[58][4] ), .D(\img_buff[59][4] ), .S0(n5077), .S1(n5061), .Y(
        n4976) );
  MX4X1 U9068 ( .A(\img_buff[60][4] ), .B(\img_buff[61][4] ), .C(
        \img_buff[62][4] ), .D(\img_buff[63][4] ), .S0(n5077), .S1(n5060), .Y(
        n4975) );
  MX4X1 U9069 ( .A(\img_buff[48][6] ), .B(\img_buff[49][6] ), .C(
        \img_buff[50][6] ), .D(\img_buff[51][6] ), .S0(n5079), .S1(n4631), .Y(
        n5018) );
  MX4X1 U9070 ( .A(\img_buff[56][6] ), .B(\img_buff[57][6] ), .C(
        \img_buff[58][6] ), .D(\img_buff[59][6] ), .S0(n5079), .S1(n4762), .Y(
        n5016) );
  MX4X1 U9071 ( .A(\img_buff[44][0] ), .B(\img_buff[45][0] ), .C(
        \img_buff[46][0] ), .D(\img_buff[47][0] ), .S0(n5624), .S1(n5639), .Y(
        n5469) );
  MX4X1 U9072 ( .A(\img_buff[28][0] ), .B(\img_buff[29][0] ), .C(
        \img_buff[30][0] ), .D(\img_buff[31][0] ), .S0(n5073), .S1(n5059), .Y(
        n4905) );
  MX4X1 U9073 ( .A(\img_buff[60][0] ), .B(\img_buff[61][0] ), .C(
        \img_buff[62][0] ), .D(\img_buff[63][0] ), .S0(n5073), .S1(n5056), .Y(
        n4895) );
  MX4X1 U9074 ( .A(\img_buff[60][0] ), .B(\img_buff[61][0] ), .C(
        \img_buff[62][0] ), .D(\img_buff[63][0] ), .S0(n4653), .S1(n5641), .Y(
        n5083) );
  MX4X1 U9075 ( .A(\img_buff[44][0] ), .B(\img_buff[45][0] ), .C(
        \img_buff[46][0] ), .D(\img_buff[47][0] ), .S0(n4653), .S1(n5642), .Y(
        n5088) );
  MX4X1 U9076 ( .A(n4903), .B(n4901), .C(n4902), .D(n4900), .S0(n5067), .S1(
        n5065), .Y(n4904) );
  MX4X1 U9077 ( .A(\img_buff[44][0] ), .B(\img_buff[45][0] ), .C(
        \img_buff[46][0] ), .D(\img_buff[47][0] ), .S0(n5073), .S1(n4631), .Y(
        n4900) );
  MX4X1 U9078 ( .A(\img_buff[36][0] ), .B(\img_buff[37][0] ), .C(
        \img_buff[38][0] ), .D(\img_buff[39][0] ), .S0(n5073), .S1(n4631), .Y(
        n4902) );
  MX4X1 U9079 ( .A(\img_buff[40][0] ), .B(\img_buff[41][0] ), .C(
        \img_buff[42][0] ), .D(\img_buff[43][0] ), .S0(n5073), .S1(n4632), .Y(
        n4901) );
  MX4X1 U9080 ( .A(\img_buff[8][2] ), .B(\img_buff[9][2] ), .C(
        \img_buff[10][2] ), .D(\img_buff[11][2] ), .S0(n5629), .S1(n5256), .Y(
        n5520) );
  MX4X1 U9081 ( .A(\img_buff[8][4] ), .B(\img_buff[9][4] ), .C(
        \img_buff[10][4] ), .D(\img_buff[11][4] ), .S0(n5632), .S1(n5644), .Y(
        n5560) );
  MX4X1 U9082 ( .A(n5512), .B(n5510), .C(n5511), .D(n5509), .S0(n5648), .S1(
        n5647), .Y(n5513) );
  MX4X1 U9083 ( .A(\img_buff[32][2] ), .B(\img_buff[33][2] ), .C(
        \img_buff[34][2] ), .D(\img_buff[35][2] ), .S0(n5629), .S1(n5266), .Y(
        n5512) );
  MX4X1 U9084 ( .A(\img_buff[40][2] ), .B(\img_buff[41][2] ), .C(
        \img_buff[42][2] ), .D(\img_buff[43][2] ), .S0(n5629), .S1(n5256), .Y(
        n5510) );
  MX4X1 U9085 ( .A(\img_buff[40][2] ), .B(\img_buff[41][2] ), .C(
        \img_buff[42][2] ), .D(\img_buff[43][2] ), .S0(n5250), .S1(n5259), .Y(
        n5129) );
  MX4X1 U9086 ( .A(\img_buff[8][2] ), .B(\img_buff[9][2] ), .C(
        \img_buff[10][2] ), .D(\img_buff[11][2] ), .S0(n5250), .S1(n5259), .Y(
        n5139) );
  MX4X1 U9087 ( .A(\img_buff[40][3] ), .B(\img_buff[41][3] ), .C(
        \img_buff[42][3] ), .D(\img_buff[43][3] ), .S0(n5436), .S1(n5450), .Y(
        n5339) );
  MX4X1 U9088 ( .A(\img_buff[8][3] ), .B(\img_buff[9][3] ), .C(
        \img_buff[10][3] ), .D(\img_buff[11][3] ), .S0(n5436), .S1(n5450), .Y(
        n5349) );
  MX4X1 U9089 ( .A(n5552), .B(n5550), .C(n5551), .D(n5549), .S0(n5648), .S1(
        n5269), .Y(n5553) );
  MX4X1 U9090 ( .A(\img_buff[40][4] ), .B(\img_buff[41][4] ), .C(
        \img_buff[42][4] ), .D(\img_buff[43][4] ), .S0(n5073), .S1(n4699), .Y(
        n5359) );
  MX4X1 U9091 ( .A(\img_buff[8][4] ), .B(\img_buff[9][4] ), .C(
        \img_buff[10][4] ), .D(\img_buff[11][4] ), .S0(n5437), .S1(n5451), .Y(
        n5369) );
  MX4X1 U9092 ( .A(\img_buff[40][4] ), .B(\img_buff[41][4] ), .C(
        \img_buff[42][4] ), .D(\img_buff[43][4] ), .S0(n5077), .S1(n5064), .Y(
        n4981) );
  MX4X1 U9093 ( .A(\img_buff[8][4] ), .B(\img_buff[9][4] ), .C(
        \img_buff[10][4] ), .D(\img_buff[11][4] ), .S0(n5078), .S1(n4695), .Y(
        n4991) );
  MX4X1 U9094 ( .A(\img_buff[8][5] ), .B(\img_buff[9][5] ), .C(
        \img_buff[10][5] ), .D(\img_buff[11][5] ), .S0(n5438), .S1(n5452), .Y(
        n5389) );
  MX4X1 U9095 ( .A(\img_buff[40][6] ), .B(\img_buff[41][6] ), .C(
        \img_buff[42][6] ), .D(\img_buff[43][6] ), .S0(n5438), .S1(n5452), .Y(
        n5399) );
  MX4X1 U9096 ( .A(\img_buff[8][6] ), .B(\img_buff[9][6] ), .C(
        \img_buff[10][6] ), .D(\img_buff[11][6] ), .S0(n5439), .S1(n5453), .Y(
        n5409) );
  MX4X1 U9097 ( .A(\img_buff[44][3] ), .B(\img_buff[45][3] ), .C(
        \img_buff[46][3] ), .D(\img_buff[47][3] ), .S0(n5076), .S1(n4695), .Y(
        n4960) );
  MX4X1 U9098 ( .A(\img_buff[36][3] ), .B(\img_buff[37][3] ), .C(
        \img_buff[38][3] ), .D(\img_buff[39][3] ), .S0(n5076), .S1(n5970), .Y(
        n4962) );
  MX4X1 U9099 ( .A(\img_buff[40][3] ), .B(\img_buff[41][3] ), .C(
        \img_buff[42][3] ), .D(\img_buff[43][3] ), .S0(n5076), .S1(n5059), .Y(
        n4961) );
  MX4X1 U9100 ( .A(\img_buff[44][7] ), .B(\img_buff[45][7] ), .C(
        \img_buff[46][7] ), .D(\img_buff[47][7] ), .S0(n5440), .S1(n5454), .Y(
        n5418) );
  MX4X1 U9101 ( .A(\img_buff[36][7] ), .B(\img_buff[37][7] ), .C(
        \img_buff[38][7] ), .D(\img_buff[39][7] ), .S0(n5440), .S1(n5454), .Y(
        n5420) );
  MX4X1 U9102 ( .A(\img_buff[40][7] ), .B(\img_buff[41][7] ), .C(
        \img_buff[42][7] ), .D(\img_buff[43][7] ), .S0(n5440), .S1(n5454), .Y(
        n5419) );
  MX4X1 U9103 ( .A(\img_buff[40][0] ), .B(\img_buff[41][0] ), .C(
        \img_buff[42][0] ), .D(\img_buff[43][0] ), .S0(n5243), .S1(n5639), .Y(
        n5470) );
  MX4X1 U9104 ( .A(\img_buff[24][0] ), .B(\img_buff[25][0] ), .C(
        \img_buff[26][0] ), .D(\img_buff[27][0] ), .S0(n5073), .S1(n5058), .Y(
        n4906) );
  MX4X1 U9105 ( .A(\img_buff[56][0] ), .B(\img_buff[57][0] ), .C(
        \img_buff[58][0] ), .D(\img_buff[59][0] ), .S0(n5073), .S1(n5062), .Y(
        n4896) );
  MX4X1 U9106 ( .A(\img_buff[56][0] ), .B(\img_buff[57][0] ), .C(
        \img_buff[58][0] ), .D(\img_buff[59][0] ), .S0(n4653), .S1(n5266), .Y(
        n5084) );
  MX4X1 U9107 ( .A(\img_buff[40][0] ), .B(\img_buff[41][0] ), .C(
        \img_buff[42][0] ), .D(\img_buff[43][0] ), .S0(n4653), .S1(n5266), .Y(
        n5089) );
  NAND4X2 U9108 ( .A(n5667), .B(n6674), .C(n6664), .D(n6659), .Y(n1820) );
  NAND4X2 U9109 ( .A(n5667), .B(n6673), .C(n6674), .D(n6659), .Y(n2454) );
  NAND4X2 U9110 ( .A(n5667), .B(n6673), .C(n6663), .D(n6659), .Y(n2137) );
  NAND4X2 U9111 ( .A(n5667), .B(n6672), .C(n6673), .D(n6663), .Y(n3405) );
  NAND4X2 U9112 ( .A(n5667), .B(n6672), .C(n6674), .D(n6664), .Y(n3088) );
  NAND4X2 U9113 ( .A(n5667), .B(n6672), .C(n6663), .D(n6664), .Y(n2771) );
  MX4X1 U9114 ( .A(\img_buff[52][3] ), .B(\img_buff[53][3] ), .C(
        \img_buff[54][3] ), .D(\img_buff[55][3] ), .S0(n5630), .S1(n5642), .Y(
        n5526) );
  MX4X1 U9115 ( .A(n5537), .B(n5535), .C(n5536), .D(n5534), .S0(n5648), .S1(
        n5647), .Y(n5538) );
  MX4X1 U9116 ( .A(\img_buff[28][3] ), .B(\img_buff[29][3] ), .C(
        \img_buff[30][3] ), .D(\img_buff[31][3] ), .S0(n5630), .S1(n5642), .Y(
        n5534) );
  MX4X1 U9117 ( .A(\img_buff[20][3] ), .B(\img_buff[21][3] ), .C(
        \img_buff[22][3] ), .D(\img_buff[23][3] ), .S0(n5630), .S1(n5642), .Y(
        n5536) );
  MX4X1 U9118 ( .A(\img_buff[24][3] ), .B(\img_buff[25][3] ), .C(
        \img_buff[26][3] ), .D(\img_buff[27][3] ), .S0(n5630), .S1(n5642), .Y(
        n5535) );
  MX4X1 U9119 ( .A(\img_buff[20][6] ), .B(\img_buff[21][6] ), .C(
        \img_buff[22][6] ), .D(\img_buff[23][6] ), .S0(n5634), .S1(n5646), .Y(
        n5596) );
  MX4X1 U9120 ( .A(\img_buff[52][6] ), .B(\img_buff[53][6] ), .C(
        \img_buff[54][6] ), .D(\img_buff[55][6] ), .S0(n5633), .S1(n5645), .Y(
        n5586) );
  MX4X1 U9121 ( .A(\img_buff[36][6] ), .B(\img_buff[37][6] ), .C(
        \img_buff[38][6] ), .D(\img_buff[39][6] ), .S0(n5634), .S1(n5646), .Y(
        n5591) );
  MX4X1 U9122 ( .A(\img_buff[4][6] ), .B(\img_buff[5][6] ), .C(
        \img_buff[6][6] ), .D(\img_buff[7][6] ), .S0(n5634), .S1(n5646), .Y(
        n5601) );
  MX4X1 U9123 ( .A(n5597), .B(n5595), .C(n5596), .D(n5594), .S0(n5650), .S1(
        n5268), .Y(n5598) );
  MX4X1 U9124 ( .A(\img_buff[16][6] ), .B(\img_buff[17][6] ), .C(
        \img_buff[18][6] ), .D(\img_buff[19][6] ), .S0(n5634), .S1(n5646), .Y(
        n5597) );
  MX4X1 U9125 ( .A(\img_buff[24][6] ), .B(\img_buff[25][6] ), .C(
        \img_buff[26][6] ), .D(\img_buff[27][6] ), .S0(n5634), .S1(n5646), .Y(
        n5595) );
  MX4X1 U9126 ( .A(\img_buff[28][6] ), .B(\img_buff[29][6] ), .C(
        \img_buff[30][6] ), .D(\img_buff[31][6] ), .S0(n5634), .S1(n5646), .Y(
        n5594) );
  MX4X1 U9127 ( .A(\img_buff[20][5] ), .B(\img_buff[21][5] ), .C(
        \img_buff[22][5] ), .D(\img_buff[23][5] ), .S0(n5633), .S1(n5645), .Y(
        n5576) );
  MX4X1 U9128 ( .A(\img_buff[4][5] ), .B(\img_buff[5][5] ), .C(
        \img_buff[6][5] ), .D(\img_buff[7][5] ), .S0(n5633), .S1(n5645), .Y(
        n5581) );
  MX4X1 U9129 ( .A(\img_buff[20][3] ), .B(\img_buff[21][3] ), .C(
        \img_buff[22][3] ), .D(\img_buff[23][3] ), .S0(n5076), .S1(n5062), .Y(
        n4967) );
  MX4X1 U9130 ( .A(\img_buff[52][3] ), .B(\img_buff[53][3] ), .C(
        \img_buff[54][3] ), .D(\img_buff[55][3] ), .S0(n5076), .S1(n5063), .Y(
        n4957) );
  MX4X1 U9131 ( .A(\img_buff[20][3] ), .B(\img_buff[21][3] ), .C(
        \img_buff[22][3] ), .D(\img_buff[23][3] ), .S0(n5629), .S1(n5260), .Y(
        n5155) );
  MX4X1 U9132 ( .A(\img_buff[52][3] ), .B(\img_buff[53][3] ), .C(
        \img_buff[54][3] ), .D(\img_buff[55][3] ), .S0(n4653), .S1(n5260), .Y(
        n5145) );
  MX4X1 U9133 ( .A(\img_buff[36][3] ), .B(\img_buff[37][3] ), .C(
        \img_buff[38][3] ), .D(\img_buff[39][3] ), .S0(n5629), .S1(n5260), .Y(
        n5150) );
  MX4X1 U9134 ( .A(\img_buff[4][3] ), .B(\img_buff[5][3] ), .C(
        \img_buff[6][3] ), .D(\img_buff[7][3] ), .S0(n5250), .S1(n5260), .Y(
        n5160) );
  MX4X1 U9135 ( .A(\img_buff[20][4] ), .B(\img_buff[21][4] ), .C(
        \img_buff[22][4] ), .D(\img_buff[23][4] ), .S0(n5251), .S1(n5261), .Y(
        n5175) );
  MX4X1 U9136 ( .A(\img_buff[52][4] ), .B(\img_buff[53][4] ), .C(
        \img_buff[54][4] ), .D(\img_buff[55][4] ), .S0(n5251), .S1(n5261), .Y(
        n5165) );
  MX4X1 U9137 ( .A(\img_buff[36][4] ), .B(\img_buff[37][4] ), .C(
        \img_buff[38][4] ), .D(\img_buff[39][4] ), .S0(n5251), .S1(n5261), .Y(
        n5170) );
  MX4X1 U9138 ( .A(\img_buff[4][4] ), .B(\img_buff[5][4] ), .C(
        \img_buff[6][4] ), .D(\img_buff[7][4] ), .S0(n5247), .S1(n5262), .Y(
        n5180) );
  MX4X1 U9139 ( .A(n5577), .B(n5575), .C(n5576), .D(n5574), .S0(n5648), .S1(
        n5269), .Y(n5578) );
  MX4X1 U9140 ( .A(\img_buff[16][5] ), .B(\img_buff[17][5] ), .C(
        \img_buff[18][5] ), .D(\img_buff[19][5] ), .S0(n5633), .S1(n5645), .Y(
        n5577) );
  MX4X1 U9141 ( .A(\img_buff[24][5] ), .B(\img_buff[25][5] ), .C(
        \img_buff[26][5] ), .D(\img_buff[27][5] ), .S0(n5633), .S1(n5645), .Y(
        n5575) );
  MX4X1 U9142 ( .A(\img_buff[28][5] ), .B(\img_buff[29][5] ), .C(
        \img_buff[30][5] ), .D(\img_buff[31][5] ), .S0(n5632), .S1(n5644), .Y(
        n5574) );
  MX4X1 U9143 ( .A(\img_buff[20][5] ), .B(\img_buff[21][5] ), .C(
        \img_buff[22][5] ), .D(\img_buff[23][5] ), .S0(n5079), .S1(n5060), .Y(
        n5007) );
  MX4X1 U9144 ( .A(\img_buff[20][5] ), .B(\img_buff[21][5] ), .C(
        \img_buff[22][5] ), .D(\img_buff[23][5] ), .S0(n5632), .S1(n5263), .Y(
        n5195) );
  MX4X1 U9145 ( .A(\img_buff[4][5] ), .B(\img_buff[5][5] ), .C(
        \img_buff[6][5] ), .D(\img_buff[7][5] ), .S0(n5244), .S1(n5263), .Y(
        n5200) );
  MX4X1 U9146 ( .A(\img_buff[20][7] ), .B(\img_buff[21][7] ), .C(
        \img_buff[22][7] ), .D(\img_buff[23][7] ), .S0(n5440), .S1(n5454), .Y(
        n5425) );
  MX4X1 U9147 ( .A(\img_buff[20][7] ), .B(\img_buff[21][7] ), .C(
        \img_buff[22][7] ), .D(\img_buff[23][7] ), .S0(n5081), .S1(n5059), .Y(
        n5047) );
  MX4X1 U9148 ( .A(\img_buff[20][6] ), .B(\img_buff[21][6] ), .C(
        \img_buff[22][6] ), .D(\img_buff[23][6] ), .S0(n5080), .S1(n5059), .Y(
        n5027) );
  MX4X1 U9149 ( .A(\img_buff[52][6] ), .B(\img_buff[53][6] ), .C(
        \img_buff[54][6] ), .D(\img_buff[55][6] ), .S0(n5079), .S1(n5970), .Y(
        n5017) );
  MX4X1 U9150 ( .A(\img_buff[36][6] ), .B(\img_buff[37][6] ), .C(
        \img_buff[38][6] ), .D(\img_buff[39][6] ), .S0(n5080), .S1(n5057), .Y(
        n5022) );
  MX4X1 U9151 ( .A(\img_buff[4][6] ), .B(\img_buff[5][6] ), .C(
        \img_buff[6][6] ), .D(\img_buff[7][6] ), .S0(n5080), .S1(n4695), .Y(
        n5032) );
  MX4X1 U9152 ( .A(\img_buff[20][6] ), .B(\img_buff[21][6] ), .C(
        \img_buff[22][6] ), .D(\img_buff[23][6] ), .S0(n5252), .S1(n5264), .Y(
        n5215) );
  MX4X1 U9153 ( .A(\img_buff[52][6] ), .B(\img_buff[53][6] ), .C(
        \img_buff[54][6] ), .D(\img_buff[55][6] ), .S0(n5244), .S1(n5263), .Y(
        n5205) );
  MX4X1 U9154 ( .A(n5156), .B(n5154), .C(n5155), .D(n5153), .S0(n5271), .S1(
        n5267), .Y(n5157) );
  MX4X1 U9155 ( .A(\img_buff[16][3] ), .B(\img_buff[17][3] ), .C(
        \img_buff[18][3] ), .D(\img_buff[19][3] ), .S0(n5251), .S1(n5260), .Y(
        n5156) );
  MX4X1 U9156 ( .A(\img_buff[24][3] ), .B(\img_buff[25][3] ), .C(
        \img_buff[26][3] ), .D(\img_buff[27][3] ), .S0(n5629), .S1(n5260), .Y(
        n5154) );
  MX4X1 U9157 ( .A(\img_buff[28][3] ), .B(\img_buff[29][3] ), .C(
        \img_buff[30][3] ), .D(\img_buff[31][3] ), .S0(n5632), .S1(n5260), .Y(
        n5153) );
  MX4X1 U9158 ( .A(n5176), .B(n5174), .C(n5175), .D(n5173), .S0(n5271), .S1(
        n5267), .Y(n5177) );
  MX4X1 U9159 ( .A(\img_buff[16][4] ), .B(\img_buff[17][4] ), .C(
        \img_buff[18][4] ), .D(\img_buff[19][4] ), .S0(n5251), .S1(n5261), .Y(
        n5176) );
  MX4X1 U9160 ( .A(\img_buff[24][4] ), .B(\img_buff[25][4] ), .C(
        \img_buff[26][4] ), .D(\img_buff[27][4] ), .S0(n5251), .S1(n5261), .Y(
        n5174) );
  MX4X1 U9161 ( .A(\img_buff[28][4] ), .B(\img_buff[29][4] ), .C(
        \img_buff[30][4] ), .D(\img_buff[31][4] ), .S0(n5251), .S1(n5261), .Y(
        n5173) );
  MX4X1 U9162 ( .A(n5196), .B(n5194), .C(n5195), .D(n5193), .S0(n5271), .S1(
        n5268), .Y(n5197) );
  MX4X1 U9163 ( .A(\img_buff[16][5] ), .B(\img_buff[17][5] ), .C(
        \img_buff[18][5] ), .D(\img_buff[19][5] ), .S0(n4653), .S1(n5263), .Y(
        n5196) );
  MX4X1 U9164 ( .A(\img_buff[24][5] ), .B(\img_buff[25][5] ), .C(
        \img_buff[26][5] ), .D(\img_buff[27][5] ), .S0(n4653), .S1(n5263), .Y(
        n5194) );
  MX4X1 U9165 ( .A(\img_buff[28][5] ), .B(\img_buff[29][5] ), .C(
        \img_buff[30][5] ), .D(\img_buff[31][5] ), .S0(n5250), .S1(n5262), .Y(
        n5193) );
  MX4X1 U9166 ( .A(n5221), .B(n5219), .C(n5220), .D(n5218), .S0(n5270), .S1(
        n5268), .Y(n5222) );
  MX4X1 U9167 ( .A(\img_buff[12][6] ), .B(\img_buff[13][6] ), .C(
        \img_buff[14][6] ), .D(\img_buff[15][6] ), .S0(n5252), .S1(n5264), .Y(
        n5218) );
  MX4X1 U9168 ( .A(\img_buff[4][6] ), .B(\img_buff[5][6] ), .C(
        \img_buff[6][6] ), .D(\img_buff[7][6] ), .S0(n5252), .S1(n5264), .Y(
        n5220) );
  MX4X1 U9169 ( .A(\img_buff[8][6] ), .B(\img_buff[9][6] ), .C(
        \img_buff[10][6] ), .D(\img_buff[11][6] ), .S0(n5252), .S1(n5264), .Y(
        n5219) );
  MX4X1 U9170 ( .A(\img_buff[32][3] ), .B(\img_buff[33][3] ), .C(
        \img_buff[34][3] ), .D(\img_buff[35][3] ), .S0(n5630), .S1(n5642), .Y(
        n5532) );
  MX4X1 U9171 ( .A(\img_buff[16][3] ), .B(\img_buff[17][3] ), .C(
        \img_buff[18][3] ), .D(\img_buff[19][3] ), .S0(n5630), .S1(n5642), .Y(
        n5537) );
  MX4X1 U9172 ( .A(\img_buff[48][3] ), .B(\img_buff[49][3] ), .C(
        \img_buff[50][3] ), .D(\img_buff[51][3] ), .S0(n5630), .S1(n5642), .Y(
        n5527) );
  MX4X1 U9173 ( .A(n5542), .B(n5540), .C(n5541), .D(n5539), .S0(n5648), .S1(
        n5647), .Y(n5543) );
  MX4X1 U9174 ( .A(\img_buff[12][3] ), .B(\img_buff[13][3] ), .C(
        \img_buff[14][3] ), .D(\img_buff[15][3] ), .S0(n5630), .S1(n5642), .Y(
        n5539) );
  MX4X1 U9175 ( .A(\img_buff[4][3] ), .B(\img_buff[5][3] ), .C(
        \img_buff[6][3] ), .D(\img_buff[7][3] ), .S0(n5630), .S1(n5642), .Y(
        n5541) );
  MX4X1 U9176 ( .A(\img_buff[8][3] ), .B(\img_buff[9][3] ), .C(
        \img_buff[10][3] ), .D(\img_buff[11][3] ), .S0(n5630), .S1(n5642), .Y(
        n5540) );
  MX4X1 U9177 ( .A(\img_buff[0][6] ), .B(\img_buff[1][6] ), .C(
        \img_buff[2][6] ), .D(\img_buff[3][6] ), .S0(n5634), .S1(n5646), .Y(
        n5602) );
  MX4X1 U9178 ( .A(\img_buff[0][5] ), .B(\img_buff[1][5] ), .C(
        \img_buff[2][5] ), .D(\img_buff[3][5] ), .S0(n5633), .S1(n5645), .Y(
        n5582) );
  MX4X1 U9179 ( .A(\img_buff[16][3] ), .B(\img_buff[17][3] ), .C(
        \img_buff[18][3] ), .D(\img_buff[19][3] ), .S0(n5076), .S1(n4632), .Y(
        n4968) );
  MX4X1 U9180 ( .A(\img_buff[48][3] ), .B(\img_buff[49][3] ), .C(
        \img_buff[50][3] ), .D(\img_buff[51][3] ), .S0(n5076), .S1(n5064), .Y(
        n4958) );
  MX4X1 U9181 ( .A(\img_buff[32][3] ), .B(\img_buff[33][3] ), .C(
        \img_buff[34][3] ), .D(\img_buff[35][3] ), .S0(n5629), .S1(n5260), .Y(
        n5151) );
  MX4X1 U9182 ( .A(\img_buff[0][3] ), .B(\img_buff[1][3] ), .C(
        \img_buff[2][3] ), .D(\img_buff[3][3] ), .S0(n5251), .S1(n5261), .Y(
        n5161) );
  MX4X1 U9183 ( .A(\img_buff[32][4] ), .B(\img_buff[33][4] ), .C(
        \img_buff[34][4] ), .D(\img_buff[35][4] ), .S0(n5251), .S1(n5261), .Y(
        n5171) );
  MX4X1 U9184 ( .A(\img_buff[0][4] ), .B(\img_buff[1][4] ), .C(
        \img_buff[2][4] ), .D(\img_buff[3][4] ), .S0(n5247), .S1(n5262), .Y(
        n5181) );
  MX4X1 U9185 ( .A(\img_buff[0][5] ), .B(\img_buff[1][5] ), .C(
        \img_buff[2][5] ), .D(\img_buff[3][5] ), .S0(n5079), .S1(n5056), .Y(
        n5013) );
  MX4X1 U9186 ( .A(\img_buff[16][5] ), .B(\img_buff[17][5] ), .C(
        \img_buff[18][5] ), .D(\img_buff[19][5] ), .S0(n5079), .S1(n4632), .Y(
        n5008) );
  MX4X1 U9187 ( .A(\img_buff[0][5] ), .B(\img_buff[1][5] ), .C(
        \img_buff[2][5] ), .D(\img_buff[3][5] ), .S0(n5632), .S1(n5263), .Y(
        n5201) );
  MX4X1 U9188 ( .A(\img_buff[0][7] ), .B(\img_buff[1][7] ), .C(
        \img_buff[2][7] ), .D(\img_buff[3][7] ), .S0(n5440), .S1(n5454), .Y(
        n5431) );
  MX4X1 U9189 ( .A(\img_buff[16][7] ), .B(\img_buff[17][7] ), .C(
        \img_buff[18][7] ), .D(\img_buff[19][7] ), .S0(n5440), .S1(n5454), .Y(
        n5426) );
  MX4X1 U9190 ( .A(\img_buff[48][7] ), .B(\img_buff[49][7] ), .C(
        \img_buff[50][7] ), .D(\img_buff[51][7] ), .S0(n5440), .S1(n5454), .Y(
        n5416) );
  MX4X1 U9191 ( .A(\img_buff[0][7] ), .B(\img_buff[1][7] ), .C(
        \img_buff[2][7] ), .D(\img_buff[3][7] ), .S0(n5081), .S1(n5970), .Y(
        n5053) );
  MX4X1 U9192 ( .A(\img_buff[16][7] ), .B(\img_buff[17][7] ), .C(
        \img_buff[18][7] ), .D(\img_buff[19][7] ), .S0(n5081), .S1(n5057), .Y(
        n5048) );
  MX4X1 U9193 ( .A(\img_buff[48][7] ), .B(\img_buff[49][7] ), .C(
        \img_buff[50][7] ), .D(\img_buff[51][7] ), .S0(n5081), .S1(n4631), .Y(
        n5038) );
  MX4X1 U9194 ( .A(\img_buff[32][6] ), .B(\img_buff[33][6] ), .C(
        \img_buff[34][6] ), .D(\img_buff[35][6] ), .S0(n5080), .S1(n5055), .Y(
        n5023) );
  MX4X1 U9195 ( .A(\img_buff[0][6] ), .B(\img_buff[1][6] ), .C(
        \img_buff[2][6] ), .D(\img_buff[3][6] ), .S0(n5080), .S1(n4631), .Y(
        n5033) );
  MX4X1 U9196 ( .A(\img_buff[0][6] ), .B(\img_buff[1][6] ), .C(
        \img_buff[2][6] ), .D(\img_buff[3][6] ), .S0(n5252), .S1(n5264), .Y(
        n5221) );
  MX4X1 U9197 ( .A(\img_buff[32][6] ), .B(\img_buff[33][6] ), .C(
        \img_buff[34][6] ), .D(\img_buff[35][6] ), .S0(n5252), .S1(n5264), .Y(
        n5211) );
  MX4X1 U9198 ( .A(\img_buff[16][6] ), .B(\img_buff[17][6] ), .C(
        \img_buff[18][6] ), .D(\img_buff[19][6] ), .S0(n5252), .S1(n5264), .Y(
        n5216) );
  MX4X1 U9199 ( .A(\img_buff[48][6] ), .B(\img_buff[49][6] ), .C(
        \img_buff[50][6] ), .D(\img_buff[51][6] ), .S0(n4653), .S1(n5263), .Y(
        n5206) );
  MX4X1 U9200 ( .A(\img_buff[12][5] ), .B(\img_buff[13][5] ), .C(
        \img_buff[14][5] ), .D(\img_buff[15][5] ), .S0(n5079), .S1(n4695), .Y(
        n5010) );
  MX4X1 U9201 ( .A(\img_buff[4][5] ), .B(\img_buff[5][5] ), .C(
        \img_buff[6][5] ), .D(\img_buff[7][5] ), .S0(n5079), .S1(n4762), .Y(
        n5012) );
  MX4X1 U9202 ( .A(\img_buff[8][5] ), .B(\img_buff[9][5] ), .C(
        \img_buff[10][5] ), .D(\img_buff[11][5] ), .S0(n5079), .S1(n5055), .Y(
        n5011) );
  MX4X1 U9203 ( .A(\img_buff[12][7] ), .B(\img_buff[13][7] ), .C(
        \img_buff[14][7] ), .D(\img_buff[15][7] ), .S0(n5081), .S1(n5062), .Y(
        n5050) );
  MX4X1 U9204 ( .A(\img_buff[4][7] ), .B(\img_buff[5][7] ), .C(
        \img_buff[6][7] ), .D(\img_buff[7][7] ), .S0(n5081), .S1(n4632), .Y(
        n5052) );
  MX4X1 U9205 ( .A(\img_buff[12][6] ), .B(\img_buff[13][6] ), .C(
        \img_buff[14][6] ), .D(\img_buff[15][6] ), .S0(n5634), .S1(n5646), .Y(
        n5599) );
  MX4X1 U9206 ( .A(n5587), .B(n5585), .C(n5586), .D(n5584), .S0(n5650), .S1(
        n5963), .Y(n5588) );
  MX4X1 U9207 ( .A(\img_buff[48][6] ), .B(\img_buff[49][6] ), .C(
        \img_buff[50][6] ), .D(\img_buff[51][6] ), .S0(n5633), .S1(n5645), .Y(
        n5587) );
  MX4X1 U9208 ( .A(\img_buff[56][6] ), .B(\img_buff[57][6] ), .C(
        \img_buff[58][6] ), .D(\img_buff[59][6] ), .S0(n5633), .S1(n5645), .Y(
        n5585) );
  MX4X1 U9209 ( .A(\img_buff[60][6] ), .B(\img_buff[61][6] ), .C(
        \img_buff[62][6] ), .D(\img_buff[63][6] ), .S0(n5633), .S1(n5645), .Y(
        n5584) );
  MX4X1 U9210 ( .A(\img_buff[12][5] ), .B(\img_buff[13][5] ), .C(
        \img_buff[14][5] ), .D(\img_buff[15][5] ), .S0(n5633), .S1(n5645), .Y(
        n5579) );
  MX4X1 U9211 ( .A(\img_buff[28][3] ), .B(\img_buff[29][3] ), .C(
        \img_buff[30][3] ), .D(\img_buff[31][3] ), .S0(n5076), .S1(n5060), .Y(
        n4965) );
  MX4X1 U9212 ( .A(\img_buff[44][3] ), .B(\img_buff[45][3] ), .C(
        \img_buff[46][3] ), .D(\img_buff[47][3] ), .S0(n5250), .S1(n5260), .Y(
        n5148) );
  MX4X1 U9213 ( .A(\img_buff[12][3] ), .B(\img_buff[13][3] ), .C(
        \img_buff[14][3] ), .D(\img_buff[15][3] ), .S0(n5629), .S1(n5260), .Y(
        n5158) );
  MX4X1 U9214 ( .A(\img_buff[44][4] ), .B(\img_buff[45][4] ), .C(
        \img_buff[46][4] ), .D(\img_buff[47][4] ), .S0(n5251), .S1(n5261), .Y(
        n5168) );
  MX4X1 U9215 ( .A(\img_buff[12][4] ), .B(\img_buff[13][4] ), .C(
        \img_buff[14][4] ), .D(\img_buff[15][4] ), .S0(n4653), .S1(n5262), .Y(
        n5178) );
  MX4X1 U9216 ( .A(\img_buff[12][5] ), .B(\img_buff[13][5] ), .C(
        \img_buff[14][5] ), .D(\img_buff[15][5] ), .S0(n5245), .S1(n5263), .Y(
        n5198) );
  MX4X1 U9217 ( .A(\img_buff[28][7] ), .B(\img_buff[29][7] ), .C(
        \img_buff[30][7] ), .D(\img_buff[31][7] ), .S0(n5440), .S1(n5454), .Y(
        n5423) );
  MX4X1 U9218 ( .A(\img_buff[28][7] ), .B(\img_buff[29][7] ), .C(
        \img_buff[30][7] ), .D(\img_buff[31][7] ), .S0(n5081), .S1(n5064), .Y(
        n5045) );
  MX4X1 U9219 ( .A(\img_buff[44][6] ), .B(\img_buff[45][6] ), .C(
        \img_buff[46][6] ), .D(\img_buff[47][6] ), .S0(n5079), .S1(n5058), .Y(
        n5020) );
  MX4X1 U9220 ( .A(\img_buff[12][6] ), .B(\img_buff[13][6] ), .C(
        \img_buff[14][6] ), .D(\img_buff[15][6] ), .S0(n5080), .S1(n5061), .Y(
        n5030) );
  MX4X1 U9221 ( .A(\img_buff[28][6] ), .B(\img_buff[29][6] ), .C(
        \img_buff[30][6] ), .D(\img_buff[31][6] ), .S0(n5252), .S1(n5264), .Y(
        n5213) );
  MX4X1 U9222 ( .A(\img_buff[60][6] ), .B(\img_buff[61][6] ), .C(
        \img_buff[62][6] ), .D(\img_buff[63][6] ), .S0(n5632), .S1(n5263), .Y(
        n5203) );
  MX4X1 U9223 ( .A(n5106), .B(n5104), .C(n5105), .D(n5103), .S0(n5272), .S1(
        n5268), .Y(n5107) );
  MX4X1 U9224 ( .A(n5146), .B(n5144), .C(n5145), .D(n5143), .S0(n5272), .S1(
        n5267), .Y(n5147) );
  MX4X1 U9225 ( .A(\img_buff[48][3] ), .B(\img_buff[49][3] ), .C(
        \img_buff[50][3] ), .D(\img_buff[51][3] ), .S0(n4653), .S1(n5260), .Y(
        n5146) );
  MX4X1 U9226 ( .A(n5166), .B(n5164), .C(n5165), .D(n5163), .S0(n5271), .S1(
        n5267), .Y(n5167) );
  MX4X1 U9227 ( .A(\img_buff[48][4] ), .B(\img_buff[49][4] ), .C(
        \img_buff[50][4] ), .D(\img_buff[51][4] ), .S0(n5251), .S1(n5261), .Y(
        n5166) );
  MX4X1 U9228 ( .A(\img_buff[56][4] ), .B(\img_buff[57][4] ), .C(
        \img_buff[58][4] ), .D(\img_buff[59][4] ), .S0(n5251), .S1(n5261), .Y(
        n5164) );
  MX4X1 U9229 ( .A(\img_buff[60][4] ), .B(\img_buff[61][4] ), .C(
        \img_buff[62][4] ), .D(\img_buff[63][4] ), .S0(n5251), .S1(n5261), .Y(
        n5163) );
  MX4X1 U9230 ( .A(n5186), .B(n5184), .C(n5185), .D(n5183), .S0(n5271), .S1(
        n5268), .Y(n5187) );
  MX4X1 U9231 ( .A(\img_buff[48][5] ), .B(\img_buff[49][5] ), .C(
        \img_buff[50][5] ), .D(\img_buff[51][5] ), .S0(n5244), .S1(n5262), .Y(
        n5186) );
  MX4X1 U9232 ( .A(\img_buff[56][5] ), .B(\img_buff[57][5] ), .C(
        \img_buff[58][5] ), .D(\img_buff[59][5] ), .S0(n5247), .S1(n5262), .Y(
        n5184) );
  MX4X1 U9233 ( .A(\img_buff[60][5] ), .B(\img_buff[61][5] ), .C(
        \img_buff[62][5] ), .D(\img_buff[63][5] ), .S0(n5632), .S1(n5262), .Y(
        n5183) );
  MX4X1 U9234 ( .A(n5532), .B(n5530), .C(n5531), .D(n5529), .S0(n5648), .S1(
        n5269), .Y(n5533) );
  MX4X1 U9235 ( .A(\img_buff[44][3] ), .B(\img_buff[45][3] ), .C(
        \img_buff[46][3] ), .D(\img_buff[47][3] ), .S0(n5630), .S1(n5642), .Y(
        n5529) );
  MX4X1 U9236 ( .A(\img_buff[36][3] ), .B(\img_buff[37][3] ), .C(
        \img_buff[38][3] ), .D(\img_buff[39][3] ), .S0(n5630), .S1(n5642), .Y(
        n5531) );
  MX4X1 U9237 ( .A(\img_buff[40][3] ), .B(\img_buff[41][3] ), .C(
        \img_buff[42][3] ), .D(\img_buff[43][3] ), .S0(n5630), .S1(n5642), .Y(
        n5530) );
  MX4X1 U9238 ( .A(\img_buff[8][6] ), .B(\img_buff[9][6] ), .C(
        \img_buff[10][6] ), .D(\img_buff[11][6] ), .S0(n5634), .S1(n5646), .Y(
        n5600) );
  MX4X1 U9239 ( .A(n5592), .B(n5590), .C(n5591), .D(n5589), .S0(n5649), .S1(
        n5963), .Y(n5593) );
  MX4X1 U9240 ( .A(\img_buff[32][6] ), .B(\img_buff[33][6] ), .C(
        \img_buff[34][6] ), .D(\img_buff[35][6] ), .S0(n5634), .S1(n5646), .Y(
        n5592) );
  MX4X1 U9241 ( .A(\img_buff[40][6] ), .B(\img_buff[41][6] ), .C(
        \img_buff[42][6] ), .D(\img_buff[43][6] ), .S0(n5633), .S1(n5645), .Y(
        n5590) );
  MX4X1 U9242 ( .A(\img_buff[44][6] ), .B(\img_buff[45][6] ), .C(
        \img_buff[46][6] ), .D(\img_buff[47][6] ), .S0(n5633), .S1(n5645), .Y(
        n5589) );
  MX4X1 U9243 ( .A(\img_buff[8][5] ), .B(\img_buff[9][5] ), .C(
        \img_buff[10][5] ), .D(\img_buff[11][5] ), .S0(n5633), .S1(n5645), .Y(
        n5580) );
  MX4X1 U9244 ( .A(\img_buff[24][3] ), .B(\img_buff[25][3] ), .C(
        \img_buff[26][3] ), .D(\img_buff[27][3] ), .S0(n5076), .S1(n5058), .Y(
        n4966) );
  MX4X1 U9245 ( .A(\img_buff[40][3] ), .B(\img_buff[41][3] ), .C(
        \img_buff[42][3] ), .D(\img_buff[43][3] ), .S0(n5250), .S1(n5260), .Y(
        n5149) );
  MX4X1 U9246 ( .A(\img_buff[8][3] ), .B(\img_buff[9][3] ), .C(
        \img_buff[10][3] ), .D(\img_buff[11][3] ), .S0(n5629), .S1(n5260), .Y(
        n5159) );
  MX4X1 U9247 ( .A(\img_buff[40][4] ), .B(\img_buff[41][4] ), .C(
        \img_buff[42][4] ), .D(\img_buff[43][4] ), .S0(n5251), .S1(n5261), .Y(
        n5169) );
  MX4X1 U9248 ( .A(\img_buff[8][4] ), .B(\img_buff[9][4] ), .C(
        \img_buff[10][4] ), .D(\img_buff[11][4] ), .S0(n5247), .S1(n5262), .Y(
        n5179) );
  MX4X1 U9249 ( .A(\img_buff[24][5] ), .B(\img_buff[25][5] ), .C(
        \img_buff[26][5] ), .D(\img_buff[27][5] ), .S0(n5079), .S1(n5064), .Y(
        n5006) );
  MX4X1 U9250 ( .A(\img_buff[8][5] ), .B(\img_buff[9][5] ), .C(
        \img_buff[10][5] ), .D(\img_buff[11][5] ), .S0(n5244), .S1(n5263), .Y(
        n5199) );
  MX4X1 U9251 ( .A(\img_buff[24][7] ), .B(\img_buff[25][7] ), .C(
        \img_buff[26][7] ), .D(\img_buff[27][7] ), .S0(n5440), .S1(n5454), .Y(
        n5424) );
  MX4X1 U9252 ( .A(\img_buff[24][7] ), .B(\img_buff[25][7] ), .C(
        \img_buff[26][7] ), .D(\img_buff[27][7] ), .S0(n5081), .S1(n5062), .Y(
        n5046) );
  MX4X1 U9253 ( .A(\img_buff[40][6] ), .B(\img_buff[41][6] ), .C(
        \img_buff[42][6] ), .D(\img_buff[43][6] ), .S0(n5079), .S1(n5061), .Y(
        n5021) );
  MX4X1 U9254 ( .A(\img_buff[8][6] ), .B(\img_buff[9][6] ), .C(
        \img_buff[10][6] ), .D(\img_buff[11][6] ), .S0(n5080), .S1(n5059), .Y(
        n5031) );
  MX4X1 U9255 ( .A(\img_buff[24][6] ), .B(\img_buff[25][6] ), .C(
        \img_buff[26][6] ), .D(\img_buff[27][6] ), .S0(n5252), .S1(n5264), .Y(
        n5214) );
  MX4X1 U9256 ( .A(\img_buff[56][6] ), .B(\img_buff[57][6] ), .C(
        \img_buff[58][6] ), .D(\img_buff[59][6] ), .S0(n5251), .S1(n5263), .Y(
        n5204) );
  MX4X1 U9257 ( .A(\img_buff[44][7] ), .B(\img_buff[45][7] ), .C(
        \img_buff[46][7] ), .D(\img_buff[47][7] ), .S0(n5081), .S1(n4632), .Y(
        n5040) );
  MX4X1 U9258 ( .A(\img_buff[36][7] ), .B(\img_buff[37][7] ), .C(
        \img_buff[38][7] ), .D(\img_buff[39][7] ), .S0(n5081), .S1(n5057), .Y(
        n5042) );
  MX4X1 U9259 ( .A(n5211), .B(n5209), .C(n5210), .D(n5208), .S0(n5271), .S1(
        n5268), .Y(n5212) );
  MX4X1 U9260 ( .A(\img_buff[44][6] ), .B(\img_buff[45][6] ), .C(
        \img_buff[46][6] ), .D(\img_buff[47][6] ), .S0(n5251), .S1(n5263), .Y(
        n5208) );
  MX4X1 U9261 ( .A(\img_buff[36][6] ), .B(\img_buff[37][6] ), .C(
        \img_buff[38][6] ), .D(\img_buff[39][6] ), .S0(n5252), .S1(n5264), .Y(
        n5210) );
  MX4X1 U9262 ( .A(\img_buff[40][6] ), .B(\img_buff[41][6] ), .C(
        \img_buff[42][6] ), .D(\img_buff[43][6] ), .S0(n5245), .S1(n5263), .Y(
        n5209) );
  OAI21X1 U9263 ( .A0(n974), .A1(n93), .B0(n6642), .Y(n4080) );
  CLKINVX1 U9264 ( .A(n4075), .Y(n6643) );
  AOI31X1 U9265 ( .A0(n4073), .A1(n5964), .A2(n6647), .B0(n944), .Y(n4076) );
  CLKINVX1 U9266 ( .A(n4067), .Y(n6647) );
  OAI211X1 U9267 ( .A0(n969), .A1(n93), .B0(n970), .C0(n6642), .Y(n968) );
  NOR4BX1 U9268 ( .AN(n5668), .B(n973), .C(n966), .D(n6649), .Y(n969) );
  OAI21XL U9269 ( .A0(n971), .A1(cmd_valid), .B0(n93), .Y(n970) );
  NAND3X1 U9270 ( .A(n974), .B(n975), .C(n5913), .Y(n973) );
  OAI2BB2XL U9271 ( .B0(n4094), .B1(n6654), .A0N(n6654), .A1N(n4095), .Y(n4625) );
  OAI2BB2XL U9272 ( .B0(n4094), .B1(n6653), .A0N(N3455), .A1N(n4095), .Y(n4626) );
  OAI2BB2XL U9273 ( .B0(n6660), .B1(n967), .A0N(N3380), .A1N(n4093), .Y(n4619)
         );
  OAI2BB2XL U9274 ( .B0(n6659), .B1(n967), .A0N(N3385), .A1N(n4093), .Y(n4620)
         );
  OAI31XL U9275 ( .A0(n4627), .A1(n4061), .A2(n4062), .B0(n4063), .Y(n4608) );
  NAND2XL U9276 ( .A(IRAM_valid), .B(n4062), .Y(n4063) );
  NOR2BX1 U9277 ( .AN(n1476), .B(n4627), .Y(n4062) );
  AO22XL U9278 ( .A0(IRAM_D[0]), .A1(n5671), .B0(n1068), .B1(n1419), .Y(n4103)
         );
  NAND4BX1 U9279 ( .AN(n1420), .B(n1421), .C(n1422), .D(n1423), .Y(n1419) );
  NOR4X1 U9280 ( .A(n1447), .B(n1448), .C(n1449), .D(n1450), .Y(n1421) );
  NOR4X1 U9281 ( .A(n1424), .B(n1425), .C(n1426), .D(n1427), .Y(n1423) );
  AO22XL U9282 ( .A0(IRAM_D[1]), .A1(n5671), .B0(n1068), .B1(n1378), .Y(n4102)
         );
  NAND4BX1 U9283 ( .AN(n1379), .B(n1380), .C(n1381), .D(n1382), .Y(n1378) );
  NOR4X1 U9284 ( .A(n1395), .B(n1396), .C(n1397), .D(n1398), .Y(n1380) );
  NOR4X1 U9285 ( .A(n1383), .B(n1384), .C(n1385), .D(n1386), .Y(n1382) );
  AO22XL U9286 ( .A0(IRAM_D[2]), .A1(n5671), .B0(n1068), .B1(n1337), .Y(n4101)
         );
  NAND4BX1 U9287 ( .AN(n1338), .B(n1339), .C(n1340), .D(n1341), .Y(n1337) );
  NOR4X1 U9288 ( .A(n1354), .B(n1355), .C(n1356), .D(n1357), .Y(n1339) );
  NOR4X1 U9289 ( .A(n1342), .B(n1343), .C(n1344), .D(n1345), .Y(n1341) );
  AO22XL U9290 ( .A0(IRAM_D[3]), .A1(n5671), .B0(n1068), .B1(n1296), .Y(n4100)
         );
  NAND4BX1 U9291 ( .AN(n1297), .B(n1298), .C(n1299), .D(n1300), .Y(n1296) );
  NOR4X1 U9292 ( .A(n1313), .B(n1314), .C(n1315), .D(n1316), .Y(n1298) );
  NOR4X1 U9293 ( .A(n1301), .B(n1302), .C(n1303), .D(n1304), .Y(n1300) );
  AO22XL U9294 ( .A0(IRAM_D[4]), .A1(n5671), .B0(n1068), .B1(n1255), .Y(n4099)
         );
  NAND4BX1 U9295 ( .AN(n1256), .B(n1257), .C(n1258), .D(n1259), .Y(n1255) );
  NOR4X1 U9296 ( .A(n1272), .B(n1273), .C(n1274), .D(n1275), .Y(n1257) );
  NOR4X1 U9297 ( .A(n1260), .B(n1261), .C(n1262), .D(n1263), .Y(n1259) );
  AO22XL U9298 ( .A0(IRAM_D[5]), .A1(n5671), .B0(n1068), .B1(n1214), .Y(n4098)
         );
  NAND4BX1 U9299 ( .AN(n1215), .B(n1216), .C(n1217), .D(n1218), .Y(n1214) );
  NOR4X1 U9300 ( .A(n1231), .B(n1232), .C(n1233), .D(n1234), .Y(n1216) );
  NOR4X1 U9301 ( .A(n1219), .B(n1220), .C(n1221), .D(n1222), .Y(n1218) );
  AO22XL U9302 ( .A0(IRAM_D[7]), .A1(n5671), .B0(n1068), .B1(n1069), .Y(n4096)
         );
  NAND4BX1 U9303 ( .AN(n1070), .B(n1071), .C(n1072), .D(n1073), .Y(n1069) );
  NOR4X1 U9304 ( .A(n1109), .B(n1110), .C(n1111), .D(n1112), .Y(n1071) );
  NOR4X1 U9305 ( .A(n1074), .B(n1075), .C(n1076), .D(n1077), .Y(n1073) );
  AO22XL U9306 ( .A0(IRAM_D[6]), .A1(n5671), .B0(n1068), .B1(n1173), .Y(n4097)
         );
  NAND4BX1 U9307 ( .AN(n1174), .B(n1175), .C(n1176), .D(n1177), .Y(n1173) );
  NOR4X1 U9308 ( .A(n1190), .B(n1191), .C(n1192), .D(n1193), .Y(n1175) );
  NOR4X1 U9309 ( .A(n1178), .B(n1179), .C(n1180), .D(n1181), .Y(n1177) );
  AND2X2 U9310 ( .A(n5667), .B(cmd_valid), .Y(n4883) );
  MX4X1 U9311 ( .A(n5236), .B(n5234), .C(n5235), .D(n5233), .S0(n5270), .S1(
        n5268), .Y(n5237) );
  MX4X1 U9312 ( .A(\img_buff[16][7] ), .B(\img_buff[17][7] ), .C(
        \img_buff[18][7] ), .D(\img_buff[19][7] ), .S0(n5253), .S1(n5265), .Y(
        n5236) );
  MX4X1 U9313 ( .A(\img_buff[24][7] ), .B(\img_buff[25][7] ), .C(
        \img_buff[26][7] ), .D(\img_buff[27][7] ), .S0(n5253), .S1(n5265), .Y(
        n5234) );
  MX4X1 U9314 ( .A(\img_buff[28][7] ), .B(\img_buff[29][7] ), .C(
        \img_buff[30][7] ), .D(\img_buff[31][7] ), .S0(n5253), .S1(n5265), .Y(
        n5233) );
  MX4X1 U9315 ( .A(\img_buff[28][7] ), .B(\img_buff[29][7] ), .C(
        \img_buff[30][7] ), .D(\img_buff[31][7] ), .S0(n5635), .S1(n5263), .Y(
        n5614) );
  MX4X1 U9316 ( .A(\img_buff[20][7] ), .B(\img_buff[21][7] ), .C(
        \img_buff[22][7] ), .D(\img_buff[23][7] ), .S0(n5635), .S1(n5646), .Y(
        n5616) );
  MX4X1 U9317 ( .A(\img_buff[24][7] ), .B(\img_buff[25][7] ), .C(
        \img_buff[26][7] ), .D(\img_buff[27][7] ), .S0(n5635), .S1(n5646), .Y(
        n5615) );
  MX4X1 U9318 ( .A(\img_buff[20][7] ), .B(\img_buff[21][7] ), .C(
        \img_buff[22][7] ), .D(\img_buff[23][7] ), .S0(n5253), .S1(n5265), .Y(
        n5235) );
  MX4X1 U9319 ( .A(\img_buff[36][7] ), .B(\img_buff[37][7] ), .C(
        \img_buff[38][7] ), .D(\img_buff[39][7] ), .S0(n5253), .S1(n5265), .Y(
        n5230) );
  MX4X1 U9320 ( .A(\img_buff[4][7] ), .B(\img_buff[5][7] ), .C(
        \img_buff[6][7] ), .D(\img_buff[7][7] ), .S0(n5253), .S1(n5265), .Y(
        n5240) );
  MX4X1 U9321 ( .A(\img_buff[0][7] ), .B(\img_buff[1][7] ), .C(
        \img_buff[2][7] ), .D(\img_buff[3][7] ), .S0(n5635), .S1(n5645), .Y(
        n5622) );
  MX4X1 U9322 ( .A(\img_buff[48][7] ), .B(\img_buff[49][7] ), .C(
        \img_buff[50][7] ), .D(\img_buff[51][7] ), .S0(n5635), .S1(n5643), .Y(
        n5607) );
  MX4X1 U9323 ( .A(\img_buff[12][7] ), .B(\img_buff[13][7] ), .C(
        \img_buff[14][7] ), .D(\img_buff[15][7] ), .S0(n5635), .S1(n5260), .Y(
        n5619) );
  MX4X1 U9324 ( .A(\img_buff[4][7] ), .B(\img_buff[5][7] ), .C(
        \img_buff[6][7] ), .D(\img_buff[7][7] ), .S0(n5635), .S1(n4749), .Y(
        n5621) );
  MX4X1 U9325 ( .A(\img_buff[8][7] ), .B(\img_buff[9][7] ), .C(
        \img_buff[10][7] ), .D(\img_buff[11][7] ), .S0(n5635), .S1(n5646), .Y(
        n5620) );
  MX4X1 U9326 ( .A(\img_buff[32][7] ), .B(\img_buff[33][7] ), .C(
        \img_buff[34][7] ), .D(\img_buff[35][7] ), .S0(n5253), .S1(n5265), .Y(
        n5231) );
  MX4X1 U9327 ( .A(\img_buff[0][7] ), .B(\img_buff[1][7] ), .C(
        \img_buff[2][7] ), .D(\img_buff[3][7] ), .S0(n5253), .S1(n5265), .Y(
        n5241) );
  MX4X1 U9328 ( .A(n5226), .B(n5224), .C(n5225), .D(n5223), .S0(n5270), .S1(
        n5268), .Y(n5227) );
  MX4X1 U9329 ( .A(\img_buff[48][7] ), .B(\img_buff[49][7] ), .C(
        \img_buff[50][7] ), .D(\img_buff[51][7] ), .S0(n5253), .S1(n5265), .Y(
        n5226) );
  MX4X1 U9330 ( .A(\img_buff[56][7] ), .B(\img_buff[57][7] ), .C(
        \img_buff[58][7] ), .D(\img_buff[59][7] ), .S0(n5252), .S1(n5264), .Y(
        n5224) );
  MX4X1 U9331 ( .A(\img_buff[60][7] ), .B(\img_buff[61][7] ), .C(
        \img_buff[62][7] ), .D(\img_buff[63][7] ), .S0(n5252), .S1(n5264), .Y(
        n5223) );
  MX4X1 U9332 ( .A(\img_buff[44][7] ), .B(\img_buff[45][7] ), .C(
        \img_buff[46][7] ), .D(\img_buff[47][7] ), .S0(n5253), .S1(n5265), .Y(
        n5228) );
  MX4X1 U9333 ( .A(\img_buff[12][7] ), .B(\img_buff[13][7] ), .C(
        \img_buff[14][7] ), .D(\img_buff[15][7] ), .S0(n5253), .S1(n5265), .Y(
        n5238) );
  MX4X1 U9334 ( .A(\img_buff[44][7] ), .B(\img_buff[45][7] ), .C(
        \img_buff[46][7] ), .D(\img_buff[47][7] ), .S0(n5635), .S1(n5261), .Y(
        n5609) );
  MX4X1 U9335 ( .A(\img_buff[36][7] ), .B(\img_buff[37][7] ), .C(
        \img_buff[38][7] ), .D(\img_buff[39][7] ), .S0(n5635), .S1(n5646), .Y(
        n5611) );
  MX4X1 U9336 ( .A(\img_buff[40][7] ), .B(\img_buff[41][7] ), .C(
        \img_buff[42][7] ), .D(\img_buff[43][7] ), .S0(n5635), .S1(n4749), .Y(
        n5610) );
  MX4X1 U9337 ( .A(\img_buff[40][7] ), .B(\img_buff[41][7] ), .C(
        \img_buff[42][7] ), .D(\img_buff[43][7] ), .S0(n5253), .S1(n5265), .Y(
        n5229) );
  MX4X1 U9338 ( .A(\img_buff[8][7] ), .B(\img_buff[9][7] ), .C(
        \img_buff[10][7] ), .D(\img_buff[11][7] ), .S0(n5253), .S1(n5265), .Y(
        n5239) );
  AND2X2 U9339 ( .A(IROM_Q[0]), .B(n93), .Y(n4884) );
  AND2X2 U9340 ( .A(IROM_Q[1]), .B(n93), .Y(n4885) );
  AND2X2 U9341 ( .A(IROM_Q[2]), .B(n93), .Y(n4886) );
  AND2X2 U9342 ( .A(IROM_Q[3]), .B(n93), .Y(n4887) );
  AND2X2 U9343 ( .A(IROM_Q[4]), .B(n93), .Y(n4888) );
  AND2X2 U9344 ( .A(IROM_Q[5]), .B(n93), .Y(n4889) );
  AND2X2 U9345 ( .A(IROM_Q[7]), .B(n93), .Y(n4890) );
  AND2X2 U9346 ( .A(IROM_Q[6]), .B(n93), .Y(n4891) );
  CLKBUFX3 U9347 ( .A(n1067), .Y(n5671) );
  OA21XL U9348 ( .A0(n1476), .A1(n93), .B0(n6642), .Y(n1067) );
  CLKINVX2 U9349 ( .A(n6692), .Y(n6654) );
  CLKINVX2 U9350 ( .A(n6688), .Y(n6658) );
  CLKINVX2 U9351 ( .A(n6690), .Y(n6656) );
  CLKINVX2 U9352 ( .A(n6687), .Y(n6653) );
  OAI22XL U9353 ( .A0(n4710), .A1(n269), .B0(n4719), .B1(n261), .Y(n1459) );
  OAI22XL U9354 ( .A0(n4710), .A1(n268), .B0(n4719), .B1(n260), .Y(n1406) );
  OAI22XL U9355 ( .A0(n4710), .A1(n267), .B0(n4719), .B1(n259), .Y(n1365) );
  OAI22XL U9356 ( .A0(n4710), .A1(n266), .B0(n4719), .B1(n258), .Y(n1324) );
  OAI22XL U9357 ( .A0(n4710), .A1(n265), .B0(n4719), .B1(n257), .Y(n1283) );
  OAI22XL U9358 ( .A0(n4710), .A1(n264), .B0(n4719), .B1(n256), .Y(n1242) );
  OAI22XL U9359 ( .A0(n4710), .A1(n262), .B0(n4719), .B1(n254), .Y(n1128) );
  OAI22XL U9360 ( .A0(n4710), .A1(n263), .B0(n4719), .B1(n255), .Y(n1201) );
  OAI22XL U9361 ( .A0(n4689), .A1(n621), .B0(n4706), .B1(n613), .Y(n1445) );
  OAI22XL U9362 ( .A0(n4689), .A1(n620), .B0(n4706), .B1(n612), .Y(n1394) );
  OAI22XL U9363 ( .A0(n4689), .A1(n619), .B0(n4706), .B1(n611), .Y(n1353) );
  OAI22XL U9364 ( .A0(n4689), .A1(n618), .B0(n4706), .B1(n610), .Y(n1312) );
  OAI22XL U9365 ( .A0(n4689), .A1(n617), .B0(n4706), .B1(n609), .Y(n1271) );
  OAI22XL U9366 ( .A0(n4689), .A1(n616), .B0(n4706), .B1(n608), .Y(n1230) );
  OAI22XL U9367 ( .A0(n4689), .A1(n614), .B0(n4706), .B1(n606), .Y(n1100) );
  OAI22XL U9368 ( .A0(n4689), .A1(n615), .B0(n4706), .B1(n607), .Y(n1189) );
  NOR4X1 U9369 ( .A(n1437), .B(n1438), .C(n1439), .D(n1440), .Y(n1422) );
  OAI22XL U9370 ( .A0(n1092), .A1(n669), .B0(n1093), .B1(n661), .Y(n1439) );
  OAI22XL U9371 ( .A0(n4704), .A1(n685), .B0(n1091), .B1(n677), .Y(n1440) );
  OAI222XL U9372 ( .A0(n1094), .A1(n701), .B0(n4692), .B1(n693), .C0(n1096), 
        .C1(n709), .Y(n1438) );
  NOR4X1 U9373 ( .A(n1387), .B(n1388), .C(n1389), .D(n1390), .Y(n1381) );
  OAI22XL U9374 ( .A0(n1092), .A1(n668), .B0(n1093), .B1(n660), .Y(n1389) );
  OAI22XL U9375 ( .A0(n4704), .A1(n684), .B0(n1091), .B1(n676), .Y(n1390) );
  OAI222XL U9376 ( .A0(n1094), .A1(n700), .B0(n4692), .B1(n692), .C0(n1096), 
        .C1(n708), .Y(n1388) );
  NOR4X1 U9377 ( .A(n1346), .B(n1347), .C(n1348), .D(n1349), .Y(n1340) );
  OAI22XL U9378 ( .A0(n1092), .A1(n667), .B0(n1093), .B1(n659), .Y(n1348) );
  OAI22XL U9379 ( .A0(n4704), .A1(n683), .B0(n1091), .B1(n675), .Y(n1349) );
  OAI222XL U9380 ( .A0(n1094), .A1(n699), .B0(n4692), .B1(n691), .C0(n1096), 
        .C1(n707), .Y(n1347) );
  NOR4X1 U9381 ( .A(n1305), .B(n1306), .C(n1307), .D(n1308), .Y(n1299) );
  OAI22XL U9382 ( .A0(n1092), .A1(n666), .B0(n1093), .B1(n658), .Y(n1307) );
  OAI22XL U9383 ( .A0(n4704), .A1(n682), .B0(n1091), .B1(n674), .Y(n1308) );
  OAI222XL U9384 ( .A0(n1094), .A1(n698), .B0(n4692), .B1(n690), .C0(n1096), 
        .C1(n706), .Y(n1306) );
  NOR4X1 U9385 ( .A(n1264), .B(n1265), .C(n1266), .D(n1267), .Y(n1258) );
  OAI22XL U9386 ( .A0(n1092), .A1(n665), .B0(n1093), .B1(n657), .Y(n1266) );
  OAI22XL U9387 ( .A0(n4704), .A1(n681), .B0(n1091), .B1(n673), .Y(n1267) );
  OAI222XL U9388 ( .A0(n1094), .A1(n697), .B0(n4692), .B1(n689), .C0(n1096), 
        .C1(n705), .Y(n1265) );
  NOR4X1 U9389 ( .A(n1223), .B(n1224), .C(n1225), .D(n1226), .Y(n1217) );
  OAI22XL U9390 ( .A0(n1092), .A1(n664), .B0(n1093), .B1(n656), .Y(n1225) );
  OAI22XL U9391 ( .A0(n4704), .A1(n680), .B0(n1091), .B1(n672), .Y(n1226) );
  OAI222XL U9392 ( .A0(n1094), .A1(n696), .B0(n4692), .B1(n688), .C0(n1096), 
        .C1(n704), .Y(n1224) );
  NOR4X1 U9393 ( .A(n1086), .B(n1087), .C(n1088), .D(n1089), .Y(n1072) );
  OAI22XL U9394 ( .A0(n1092), .A1(n662), .B0(n1093), .B1(n654), .Y(n1088) );
  OAI22XL U9395 ( .A0(n4704), .A1(n678), .B0(n1091), .B1(n670), .Y(n1089) );
  OAI222XL U9396 ( .A0(n1094), .A1(n694), .B0(n4692), .B1(n686), .C0(n1096), 
        .C1(n702), .Y(n1087) );
  NOR4X1 U9397 ( .A(n1182), .B(n1183), .C(n1184), .D(n1185), .Y(n1176) );
  OAI22XL U9398 ( .A0(n1092), .A1(n663), .B0(n1093), .B1(n655), .Y(n1184) );
  OAI22XL U9399 ( .A0(n4704), .A1(n679), .B0(n1091), .B1(n671), .Y(n1185) );
  OAI222XL U9400 ( .A0(n1094), .A1(n695), .B0(n4692), .B1(n687), .C0(n1096), 
        .C1(n703), .Y(n1183) );
  NOR4X1 U9401 ( .A(n1456), .B(n1457), .C(n1458), .D(n1459), .Y(n1455) );
  OAI22XL U9402 ( .A0(n4690), .A1(n221), .B0(n4717), .B1(n213), .Y(n1456) );
  OAI22XL U9403 ( .A0(n1133), .A1(n237), .B0(n1134), .B1(n229), .Y(n1457) );
  OAI22XL U9404 ( .A0(n4691), .A1(n253), .B0(n1132), .B1(n245), .Y(n1458) );
  NOR4X1 U9405 ( .A(n1403), .B(n1404), .C(n1405), .D(n1406), .Y(n1402) );
  OAI22XL U9406 ( .A0(n4690), .A1(n220), .B0(n4717), .B1(n212), .Y(n1403) );
  OAI22XL U9407 ( .A0(n1133), .A1(n236), .B0(n1134), .B1(n228), .Y(n1404) );
  OAI22XL U9408 ( .A0(n4691), .A1(n252), .B0(n1132), .B1(n244), .Y(n1405) );
  NOR4X1 U9409 ( .A(n1362), .B(n1363), .C(n1364), .D(n1365), .Y(n1361) );
  OAI22XL U9410 ( .A0(n4690), .A1(n219), .B0(n4717), .B1(n211), .Y(n1362) );
  OAI22XL U9411 ( .A0(n1133), .A1(n235), .B0(n1134), .B1(n227), .Y(n1363) );
  OAI22XL U9412 ( .A0(n4691), .A1(n251), .B0(n1132), .B1(n243), .Y(n1364) );
  NOR4X1 U9413 ( .A(n1321), .B(n1322), .C(n1323), .D(n1324), .Y(n1320) );
  OAI22XL U9414 ( .A0(n4690), .A1(n218), .B0(n4717), .B1(n210), .Y(n1321) );
  OAI22XL U9415 ( .A0(n1133), .A1(n234), .B0(n1134), .B1(n226), .Y(n1322) );
  OAI22XL U9416 ( .A0(n4691), .A1(n250), .B0(n1132), .B1(n242), .Y(n1323) );
  NOR4X1 U9417 ( .A(n1280), .B(n1281), .C(n1282), .D(n1283), .Y(n1279) );
  OAI22XL U9418 ( .A0(n4690), .A1(n217), .B0(n4717), .B1(n209), .Y(n1280) );
  OAI22XL U9419 ( .A0(n1133), .A1(n233), .B0(n1134), .B1(n225), .Y(n1281) );
  OAI22XL U9420 ( .A0(n4691), .A1(n249), .B0(n1132), .B1(n241), .Y(n1282) );
  NOR4X1 U9421 ( .A(n1239), .B(n1240), .C(n1241), .D(n1242), .Y(n1238) );
  OAI22XL U9422 ( .A0(n4690), .A1(n216), .B0(n4717), .B1(n208), .Y(n1239) );
  OAI22XL U9423 ( .A0(n1133), .A1(n232), .B0(n1134), .B1(n224), .Y(n1240) );
  OAI22XL U9424 ( .A0(n4691), .A1(n248), .B0(n1132), .B1(n240), .Y(n1241) );
  NOR4X1 U9425 ( .A(n1125), .B(n1126), .C(n1127), .D(n1128), .Y(n1124) );
  OAI22XL U9426 ( .A0(n4690), .A1(n214), .B0(n4717), .B1(n206), .Y(n1125) );
  OAI22XL U9427 ( .A0(n1133), .A1(n230), .B0(n1134), .B1(n222), .Y(n1126) );
  OAI22XL U9428 ( .A0(n4691), .A1(n246), .B0(n1132), .B1(n238), .Y(n1127) );
  NOR4X1 U9429 ( .A(n1198), .B(n1199), .C(n1200), .D(n1201), .Y(n1197) );
  OAI22XL U9430 ( .A0(n4690), .A1(n215), .B0(n4717), .B1(n207), .Y(n1198) );
  OAI22XL U9431 ( .A0(n1133), .A1(n231), .B0(n1134), .B1(n223), .Y(n1199) );
  OAI22XL U9432 ( .A0(n4691), .A1(n247), .B0(n1132), .B1(n239), .Y(n1200) );
  OAI2BB2XL U9433 ( .B0(n966), .B1(n93), .A0N(n93), .A1N(cmd_valid), .Y(
        next_state) );
  NAND2X1 U9434 ( .A(n6642), .B(n4091), .Y(n4614) );
  OAI2BB1XL U9435 ( .A0N(n93), .A1N(n971), .B0(IROM_rd), .Y(n4091) );
  OR4X1 U9436 ( .A(n1442), .B(n1443), .C(n1444), .D(n1445), .Y(n1437) );
  OAI22XL U9437 ( .A0(n4688), .A1(n637), .B0(n4703), .B1(n629), .Y(n1442) );
  OAI22XL U9438 ( .A0(n1105), .A1(n653), .B0(n1106), .B1(n645), .Y(n1443) );
  OAI22XL U9439 ( .A0(n4686), .A1(n605), .B0(n1104), .B1(n597), .Y(n1444) );
  OR4X1 U9440 ( .A(n1391), .B(n1392), .C(n1393), .D(n1394), .Y(n1387) );
  OAI22XL U9441 ( .A0(n4688), .A1(n636), .B0(n4703), .B1(n628), .Y(n1391) );
  OAI22XL U9442 ( .A0(n1105), .A1(n652), .B0(n1106), .B1(n644), .Y(n1392) );
  OAI22XL U9443 ( .A0(n4686), .A1(n604), .B0(n1104), .B1(n596), .Y(n1393) );
  OR4X1 U9444 ( .A(n1350), .B(n1351), .C(n1352), .D(n1353), .Y(n1346) );
  OAI22XL U9445 ( .A0(n4688), .A1(n635), .B0(n4703), .B1(n627), .Y(n1350) );
  OAI22XL U9446 ( .A0(n1105), .A1(n651), .B0(n1106), .B1(n643), .Y(n1351) );
  OAI22XL U9447 ( .A0(n4686), .A1(n603), .B0(n1104), .B1(n595), .Y(n1352) );
  OR4X1 U9448 ( .A(n1309), .B(n1310), .C(n1311), .D(n1312), .Y(n1305) );
  OAI22XL U9449 ( .A0(n4688), .A1(n634), .B0(n4703), .B1(n626), .Y(n1309) );
  OAI22XL U9450 ( .A0(n1105), .A1(n650), .B0(n1106), .B1(n642), .Y(n1310) );
  OAI22XL U9451 ( .A0(n4686), .A1(n602), .B0(n1104), .B1(n594), .Y(n1311) );
  OR4X1 U9452 ( .A(n1268), .B(n1269), .C(n1270), .D(n1271), .Y(n1264) );
  OAI22XL U9453 ( .A0(n4688), .A1(n633), .B0(n4703), .B1(n625), .Y(n1268) );
  OAI22XL U9454 ( .A0(n1105), .A1(n649), .B0(n1106), .B1(n641), .Y(n1269) );
  OAI22XL U9455 ( .A0(n4686), .A1(n601), .B0(n1104), .B1(n593), .Y(n1270) );
  OR4X1 U9456 ( .A(n1227), .B(n1228), .C(n1229), .D(n1230), .Y(n1223) );
  OAI22XL U9457 ( .A0(n4688), .A1(n632), .B0(n4703), .B1(n624), .Y(n1227) );
  OAI22XL U9458 ( .A0(n1105), .A1(n648), .B0(n1106), .B1(n640), .Y(n1228) );
  OAI22XL U9459 ( .A0(n4686), .A1(n600), .B0(n1104), .B1(n592), .Y(n1229) );
  OR4X1 U9460 ( .A(n1097), .B(n1098), .C(n1099), .D(n1100), .Y(n1086) );
  OAI22XL U9461 ( .A0(n4688), .A1(n630), .B0(n4703), .B1(n622), .Y(n1097) );
  OAI22XL U9462 ( .A0(n1105), .A1(n646), .B0(n1106), .B1(n638), .Y(n1098) );
  OAI22XL U9463 ( .A0(n4686), .A1(n598), .B0(n1104), .B1(n590), .Y(n1099) );
  OR4X1 U9464 ( .A(n1186), .B(n1187), .C(n1188), .D(n1189), .Y(n1182) );
  OAI22XL U9465 ( .A0(n4688), .A1(n631), .B0(n4703), .B1(n623), .Y(n1186) );
  OAI22XL U9466 ( .A0(n1105), .A1(n647), .B0(n1106), .B1(n639), .Y(n1187) );
  OAI22XL U9467 ( .A0(n4686), .A1(n599), .B0(n1104), .B1(n591), .Y(n1188) );
  NAND3X2 U9468 ( .A(n6677), .B(n6661), .C(n6675), .Y(n1687) );
  NAND3X2 U9469 ( .A(n6677), .B(n6662), .C(n6676), .Y(n1599) );
  NAND3X2 U9470 ( .A(n6676), .B(n6660), .C(n6675), .Y(n1731) );
  NAND3X2 U9471 ( .A(n6676), .B(n6677), .C(n6675), .Y(n1775) );
  CLKINVX2 U9472 ( .A(n6673), .Y(n6664) );
  CLKINVX2 U9473 ( .A(n6674), .Y(n6663) );
  CLKINVX2 U9474 ( .A(n6672), .Y(n6659) );
  NAND3X2 U9475 ( .A(n6661), .B(n6662), .C(n6677), .Y(n1511) );
  NAND3X2 U9476 ( .A(n6660), .B(n6661), .C(n6675), .Y(n1643) );
  NAND3X2 U9477 ( .A(n6660), .B(n6662), .C(n6676), .Y(n1555) );
  NOR2X1 U9478 ( .A(cmd_reg[2]), .B(cmd_reg[1]), .Y(n4057) );
  NAND3X1 U9479 ( .A(cmd_reg[0]), .B(n4057), .C(cmd_reg[3]), .Y(n1034) );
  NAND3X2 U9480 ( .A(cmd_reg[2]), .B(n4059), .C(cmd_reg[1]), .Y(n4000) );
  NOR2X1 U9481 ( .A(cmd_reg[3]), .B(cmd_reg[0]), .Y(n4060) );
  CLKBUFX3 U9482 ( .A(n972), .Y(n5668) );
  OAI32X1 U9483 ( .A0(n944), .A1(n4073), .A2(n5964), .B0(n4074), .B1(n4068), 
        .Y(n4071) );
  NAND2X1 U9484 ( .A(n944), .B(n5964), .Y(n4074) );
  CLKBUFX3 U9485 ( .A(cur_state), .Y(n5954) );
  XNOR2X4 U9486 ( .A(n5674), .B(n5955), .Y(N3327) );
  XNOR2X4 U9487 ( .A(n5674), .B(n4829), .Y(N3321) );
  MX4X2 U9488 ( .A(n5292), .B(n5282), .C(n5287), .D(n5277), .S0(N3334), .S1(
        N3333), .Y(N3367) );
  MX4X2 U9489 ( .A(n5332), .B(n5322), .C(n5327), .D(n5317), .S0(N3334), .S1(
        N3333), .Y(N3365) );
  AOI31XL U9490 ( .A0(n6335), .A1(n6321), .A2(n6320), .B0(n6332), .Y(n6323) );
  XNOR2X4 U9491 ( .A(n5674), .B(n5973), .Y(N3333) );
  AO21X1 U9492 ( .A0(n5971), .A1(n5963), .B0(n5972), .Y(N3331) );
  NOR2X1 U9493 ( .A(n5674), .B(n5973), .Y(n5974) );
  NAND2BX1 U9494 ( .AN(n5659), .B(n5653), .Y(n5997) );
  NAND2X1 U9495 ( .A(N3353), .B(n6005), .Y(n5983) );
  NAND2X1 U9496 ( .A(n4667), .B(n6004), .Y(n5993) );
  NAND2BX1 U9497 ( .AN(n5656), .B(N3357), .Y(n5978) );
  NOR2BX1 U9498 ( .AN(N3359), .B(N3351), .Y(n5976) );
  NAND2BX1 U9499 ( .AN(N3357), .B(n5656), .Y(n5988) );
  AND2X1 U9500 ( .A(n5978), .B(n5988), .Y(n5985) );
  NOR2X1 U9501 ( .A(n6004), .B(n4667), .Y(n5990) );
  NOR2BX1 U9502 ( .AN(N3355), .B(n5654), .Y(n5979) );
  NOR2BX1 U9503 ( .AN(n5654), .B(N3355), .Y(n5991) );
  NOR2BX1 U9504 ( .AN(n5659), .B(n5653), .Y(n5995) );
  AOI211X1 U9505 ( .A0(n5980), .A1(n5992), .B0(n5979), .C0(n5995), .Y(n5981)
         );
  NOR3BXL U9506 ( .AN(n5997), .B(n5996), .C(n5981), .Y(n5982) );
  AOI31X1 U9507 ( .A0(n6006), .A1(n5983), .A2(n5999), .B0(n6002), .Y(n5984) );
  NOR2BX1 U9508 ( .AN(N3351), .B(N3359), .Y(n5987) );
  AOI211X1 U9509 ( .A0(n5998), .A1(n5997), .B0(n5996), .C0(n5995), .Y(n6000)
         );
  OAI31XL U9510 ( .A0(n6002), .A1(n6001), .A2(n6000), .B0(n5999), .Y(N4817) );
  NAND2BX1 U9511 ( .AN(n5661), .B(n5653), .Y(n6030) );
  NAND2X1 U9512 ( .A(n5660), .B(n6037), .Y(n6016) );
  NAND2X1 U9513 ( .A(n5663), .B(n6067), .Y(n6026) );
  NAND2BX1 U9514 ( .AN(n5656), .B(n5664), .Y(n6011) );
  NOR2BX1 U9515 ( .AN(n5666), .B(N3351), .Y(n6009) );
  NAND2BX1 U9516 ( .AN(n5664), .B(n5656), .Y(n6021) );
  NOR2X1 U9517 ( .A(n6004), .B(n5663), .Y(n6023) );
  NOR2BX1 U9518 ( .AN(n5662), .B(n5654), .Y(n6012) );
  NOR2BX1 U9519 ( .AN(n5654), .B(n5662), .Y(n6024) );
  NOR2BX1 U9520 ( .AN(n5661), .B(n5653), .Y(n6028) );
  AOI211X1 U9521 ( .A0(n6013), .A1(n6025), .B0(n6012), .C0(n6028), .Y(n6014)
         );
  NOR3BXL U9522 ( .AN(n6030), .B(n6029), .C(n6014), .Y(n6015) );
  NAND2X1 U9523 ( .A(N3360), .B(n6007), .Y(n6032) );
  AOI31X1 U9524 ( .A0(n6038), .A1(n6016), .A2(n6032), .B0(n6035), .Y(n6017) );
  NOR2BX1 U9525 ( .AN(N3351), .B(n5666), .Y(n6020) );
  OAI2BB1X1 U9526 ( .A0N(n6020), .A1N(n5657), .B0(n5665), .Y(n6019) );
  OAI211X1 U9527 ( .A0(n5657), .A1(n6020), .B0(n6019), .C0(n6018), .Y(n6022)
         );
  NAND3BX1 U9528 ( .AN(n6023), .B(n6022), .C(n6021), .Y(n6027) );
  AOI31X1 U9529 ( .A0(n6027), .A1(n6026), .A2(n6025), .B0(n6024), .Y(n6031) );
  AOI211X1 U9530 ( .A0(n6031), .A1(n6030), .B0(n6029), .C0(n6028), .Y(n6033)
         );
  OAI31XL U9531 ( .A0(n6035), .A1(n6034), .A2(n6033), .B0(n6032), .Y(N4818) );
  NAND2BX1 U9532 ( .AN(n6064), .B(n6047), .Y(n6059) );
  NOR2BX1 U9533 ( .AN(n5457), .B(N3351), .Y(n6040) );
  AO21X1 U9534 ( .A0(n6066), .A1(n6040), .B0(n5922), .Y(n6039) );
  AND2X1 U9535 ( .A(n6042), .B(n6051), .Y(n6049) );
  OAI211X1 U9536 ( .A0(n6040), .A1(n6066), .B0(n6039), .C0(n6049), .Y(n6041)
         );
  NOR2X1 U9537 ( .A(n6067), .B(n5930), .Y(n6053) );
  AOI31X1 U9538 ( .A0(n6056), .A1(n6042), .A2(n6041), .B0(n6053), .Y(n6044) );
  NOR2X1 U9539 ( .A(n6043), .B(n6054), .Y(n6055) );
  AOI211X1 U9540 ( .A0(n6044), .A1(n6055), .B0(n6043), .C0(n6058), .Y(n6045)
         );
  AOI31X1 U9541 ( .A0(n6069), .A1(n6047), .A2(n6062), .B0(n6065), .Y(n6048) );
  AOI31X1 U9542 ( .A0(n6057), .A1(n6056), .A2(n6055), .B0(n6054), .Y(n6061) );
  AOI211X1 U9543 ( .A0(n6061), .A1(n6060), .B0(n6059), .C0(n6058), .Y(n6063)
         );
  OAI31XL U9544 ( .A0(n6065), .A1(n6064), .A2(n6063), .B0(n6062), .Y(N4819) );
  NAND2X1 U9545 ( .A(n5652), .B(n6100), .Y(n6079) );
  NAND2X1 U9546 ( .A(n5655), .B(n6099), .Y(n6089) );
  NAND2BX1 U9547 ( .AN(N3357), .B(n5656), .Y(n6074) );
  NOR2BX1 U9548 ( .AN(N3351), .B(N3359), .Y(n6072) );
  AO21X1 U9549 ( .A0(n6098), .A1(n6072), .B0(n5657), .Y(n6071) );
  NAND2BX1 U9550 ( .AN(n5656), .B(N3357), .Y(n6084) );
  OAI211X1 U9551 ( .A0(n6072), .A1(n6098), .B0(n6071), .C0(n6081), .Y(n6073)
         );
  NOR2X1 U9552 ( .A(n6099), .B(n5655), .Y(n6086) );
  AOI31X1 U9553 ( .A0(n6089), .A1(n6074), .A2(n6073), .B0(n6086), .Y(n6076) );
  NOR2BX1 U9554 ( .AN(n5654), .B(N3355), .Y(n6075) );
  NOR2BX1 U9555 ( .AN(N3355), .B(n5654), .Y(n6087) );
  AOI31X1 U9556 ( .A0(n6102), .A1(n6079), .A2(n6095), .B0(n6097), .Y(n6080) );
  NOR2BX1 U9557 ( .AN(N3359), .B(N3351), .Y(n6083) );
  NAND2BX1 U9558 ( .AN(n5661), .B(n5659), .Y(n6125) );
  NAND2X1 U9559 ( .A(n5660), .B(n6133), .Y(n6111) );
  NAND2X1 U9560 ( .A(n5663), .B(n6132), .Y(n6121) );
  NAND2BX1 U9561 ( .AN(N3357), .B(n5664), .Y(n6106) );
  NOR2BX1 U9562 ( .AN(n5666), .B(N3359), .Y(n6104) );
  AO21X1 U9563 ( .A0(n6131), .A1(n6104), .B0(n5665), .Y(n6103) );
  NAND2BX1 U9564 ( .AN(n5664), .B(N3357), .Y(n6116) );
  AND2X1 U9565 ( .A(n6106), .B(n6116), .Y(n6113) );
  OAI211X1 U9566 ( .A0(n6104), .A1(n6131), .B0(n6103), .C0(n6113), .Y(n6105)
         );
  NOR2X1 U9567 ( .A(n6132), .B(N3364), .Y(n6118) );
  AOI31X1 U9568 ( .A0(n6121), .A1(n6106), .A2(n6105), .B0(n6118), .Y(n6108) );
  NOR2BX1 U9569 ( .AN(n5662), .B(N3355), .Y(n6107) );
  NOR2BX1 U9570 ( .AN(N3355), .B(n5662), .Y(n6119) );
  NOR2BX1 U9571 ( .AN(n5661), .B(n5659), .Y(n6123) );
  AOI31X1 U9572 ( .A0(n6134), .A1(n6111), .A2(n6127), .B0(n6130), .Y(n6112) );
  NOR2BX1 U9573 ( .AN(N3359), .B(n5666), .Y(n6115) );
  OAI211X1 U9574 ( .A0(N3358), .A1(n6115), .B0(n6114), .C0(n6113), .Y(n6117)
         );
  NAND3BX1 U9575 ( .AN(n6118), .B(n6117), .C(n6116), .Y(n6122) );
  AOI31X1 U9576 ( .A0(n6122), .A1(n6121), .A2(n6120), .B0(n6119), .Y(n6126) );
  NAND2BX1 U9577 ( .AN(n6160), .B(n6143), .Y(n6155) );
  NAND2BX1 U9578 ( .AN(N3357), .B(n5926), .Y(n6138) );
  NOR2BX1 U9579 ( .AN(n5457), .B(N3359), .Y(n6136) );
  AO21X1 U9580 ( .A0(n4817), .A1(n6136), .B0(n5922), .Y(n6135) );
  OAI211X1 U9581 ( .A0(n6136), .A1(n6098), .B0(n6135), .C0(n6145), .Y(n6137)
         );
  NOR2X1 U9582 ( .A(n6162), .B(n5930), .Y(n6149) );
  AOI31X1 U9583 ( .A0(n6152), .A1(n6138), .A2(n6137), .B0(n6149), .Y(n6140) );
  NOR2BX1 U9584 ( .AN(n5936), .B(N3355), .Y(n6139) );
  NAND2X1 U9585 ( .A(n5948), .B(n6165), .Y(n6158) );
  NOR2X1 U9586 ( .A(n6165), .B(n5948), .Y(n6161) );
  AOI31X1 U9587 ( .A0(n6164), .A1(n6143), .A2(n6158), .B0(n6161), .Y(n6144) );
  OAI211X1 U9588 ( .A0(N3358), .A1(n4651), .B0(n6146), .C0(n6145), .Y(n6148)
         );
  NAND3BX1 U9589 ( .AN(n6149), .B(n6148), .C(n6147), .Y(n6153) );
  AOI31X1 U9590 ( .A0(n6153), .A1(n6152), .A2(n6151), .B0(n6150), .Y(n6157) );
  NAND2BX1 U9591 ( .AN(n5653), .B(n5661), .Y(n6188) );
  NAND2X1 U9592 ( .A(n5652), .B(n6258), .Y(n6174) );
  NAND2X1 U9593 ( .A(n5655), .B(n4654), .Y(n6184) );
  NAND2BX1 U9594 ( .AN(n5664), .B(n5656), .Y(n6169) );
  NOR2BX1 U9595 ( .AN(N3351), .B(n5666), .Y(n6167) );
  AO21X1 U9596 ( .A0(n6194), .A1(n6167), .B0(n5657), .Y(n6166) );
  NAND2BX1 U9597 ( .AN(n5656), .B(n5664), .Y(n6179) );
  AND2X1 U9598 ( .A(n6169), .B(n6179), .Y(n6176) );
  OAI211X1 U9599 ( .A0(n6167), .A1(n6194), .B0(n6166), .C0(n6176), .Y(n6168)
         );
  AOI31X1 U9600 ( .A0(n6184), .A1(n6169), .A2(n6168), .B0(n6181), .Y(n6171) );
  NOR2BX1 U9601 ( .AN(n5654), .B(n5662), .Y(n6170) );
  NOR2BX1 U9602 ( .AN(n5662), .B(n5654), .Y(n6182) );
  NOR2BX1 U9603 ( .AN(n5653), .B(n5661), .Y(n6186) );
  AOI31X1 U9604 ( .A0(n6196), .A1(n6174), .A2(n6190), .B0(n6193), .Y(n6175) );
  NOR2BX1 U9605 ( .AN(n5666), .B(N3351), .Y(n6178) );
  OAI211X1 U9606 ( .A0(n5665), .A1(n6178), .B0(n6177), .C0(n6176), .Y(n6180)
         );
  NAND3BX1 U9607 ( .AN(n6181), .B(n6180), .C(n6179), .Y(n6185) );
  AOI31X1 U9608 ( .A0(n6185), .A1(n6184), .A2(n6183), .B0(n6182), .Y(n6189) );
  AOI211X1 U9609 ( .A0(n6189), .A1(n6188), .B0(n6187), .C0(n6186), .Y(n6191)
         );
  NAND2BX1 U9610 ( .AN(n5659), .B(n5661), .Y(n6219) );
  NAND2X1 U9611 ( .A(N3353), .B(n6227), .Y(n6205) );
  NAND2BX1 U9612 ( .AN(n5664), .B(N3357), .Y(n6200) );
  NOR2BX1 U9613 ( .AN(N3359), .B(n5666), .Y(n6198) );
  AO21X1 U9614 ( .A0(n6225), .A1(n6198), .B0(N3358), .Y(n6197) );
  NAND2BX1 U9615 ( .AN(N3357), .B(n5664), .Y(n6210) );
  AND2X1 U9616 ( .A(n6200), .B(n6210), .Y(n6207) );
  OAI211X1 U9617 ( .A0(n6198), .A1(n6225), .B0(n6197), .C0(n6207), .Y(n6199)
         );
  AOI31X1 U9618 ( .A0(n6215), .A1(n6200), .A2(n6199), .B0(n6212), .Y(n6202) );
  NOR2BX1 U9619 ( .AN(N3355), .B(n5662), .Y(n6201) );
  NOR2BX1 U9620 ( .AN(n5662), .B(N3355), .Y(n6213) );
  NOR2BX1 U9621 ( .AN(n5659), .B(n5661), .Y(n6217) );
  AOI31X1 U9622 ( .A0(n6229), .A1(n6205), .A2(n6221), .B0(n6224), .Y(n6206) );
  NOR2BX1 U9623 ( .AN(n5666), .B(N3359), .Y(n6209) );
  OAI211X1 U9624 ( .A0(n5665), .A1(n6209), .B0(n6208), .C0(n6207), .Y(n6211)
         );
  NAND3BX1 U9625 ( .AN(n6212), .B(n6211), .C(n6210), .Y(n6216) );
  AOI31X1 U9626 ( .A0(n6216), .A1(n6215), .A2(n6214), .B0(n6213), .Y(n6220) );
  AOI211X1 U9627 ( .A0(n6220), .A1(n6219), .B0(n6218), .C0(n6217), .Y(n6222)
         );
  NOR2X1 U9628 ( .A(n6258), .B(n5945), .Y(n6255) );
  NAND2X1 U9629 ( .A(n5944), .B(n6258), .Y(n6238) );
  NAND2X1 U9630 ( .A(n5929), .B(n4654), .Y(n6247) );
  NAND2BX1 U9631 ( .AN(n5664), .B(n5926), .Y(n6233) );
  AO21X1 U9632 ( .A0(n6194), .A1(n6231), .B0(n5922), .Y(n6230) );
  NAND2BX1 U9633 ( .AN(n5926), .B(n5664), .Y(n6242) );
  OAI211X1 U9634 ( .A0(n6231), .A1(n6225), .B0(n6230), .C0(n6240), .Y(n6232)
         );
  NOR2X1 U9635 ( .A(n6257), .B(n5930), .Y(n6244) );
  AOI31X1 U9636 ( .A0(n6247), .A1(n6233), .A2(n6232), .B0(n6244), .Y(n6235) );
  NOR2BX1 U9637 ( .AN(n5936), .B(n5662), .Y(n6234) );
  NOR2BX1 U9638 ( .AN(n5662), .B(n5936), .Y(n6245) );
  NOR2X1 U9639 ( .A(n6234), .B(n6245), .Y(n6246) );
  AOI211X1 U9640 ( .A0(n6235), .A1(n6246), .B0(n6234), .C0(n6249), .Y(n6236)
         );
  NOR2X1 U9641 ( .A(n6260), .B(n5948), .Y(n6256) );
  OAI211X1 U9642 ( .A0(n5665), .A1(n6319), .B0(n6241), .C0(n6240), .Y(n6243)
         );
  NAND3BX1 U9643 ( .AN(n6244), .B(n6243), .C(n6242), .Y(n6248) );
  AOI31X1 U9644 ( .A0(n6248), .A1(n6247), .A2(n6246), .B0(n6245), .Y(n6252) );
  AOI211X1 U9645 ( .A0(n6252), .A1(n6251), .B0(n6250), .C0(n6249), .Y(n6254)
         );
  NAND2X1 U9646 ( .A(n5652), .B(n5946), .Y(n6269) );
  AO21X1 U9647 ( .A0(n5923), .A1(n6262), .B0(n5657), .Y(n6261) );
  OAI211X1 U9648 ( .A0(n6262), .A1(n5923), .B0(n6261), .C0(n6271), .Y(n6263)
         );
  NOR2X1 U9649 ( .A(n5931), .B(n5655), .Y(n6276) );
  AOI31X1 U9650 ( .A0(n6279), .A1(n6264), .A2(n6263), .B0(n6276), .Y(n6266) );
  NOR2BX1 U9651 ( .AN(n5654), .B(n5935), .Y(n6265) );
  NOR2BX1 U9652 ( .AN(n5936), .B(n5654), .Y(n6277) );
  NAND2X1 U9653 ( .A(n5651), .B(n5950), .Y(n6285) );
  AOI31X1 U9654 ( .A0(n6289), .A1(n6269), .A2(n6285), .B0(n6288), .Y(n6270) );
  OAI2BB1X1 U9655 ( .A0N(n6273), .A1N(n5922), .B0(n5657), .Y(n6272) );
  OAI211X1 U9656 ( .A0(n5922), .A1(n6273), .B0(n6272), .C0(n6271), .Y(n6275)
         );
  NAND3BX1 U9657 ( .AN(n6276), .B(n6275), .C(n6274), .Y(n6280) );
  AOI31X1 U9658 ( .A0(n6280), .A1(n6279), .A2(n6278), .B0(n6277), .Y(n6284) );
  AOI211X1 U9659 ( .A0(n6284), .A1(n6283), .B0(n6282), .C0(n6281), .Y(n6286)
         );
  NAND2X1 U9660 ( .A(N3353), .B(n5946), .Y(n6297) );
  NAND2BX1 U9661 ( .AN(n6315), .B(n6297), .Y(n6310) );
  AO21X1 U9662 ( .A0(n5923), .A1(n4651), .B0(N3358), .Y(n6290) );
  AND2X1 U9663 ( .A(n6293), .B(n6302), .Y(n6299) );
  OAI211X1 U9664 ( .A0(n4651), .A1(n5923), .B0(n6290), .C0(n6299), .Y(n6292)
         );
  NOR2X1 U9665 ( .A(n5932), .B(n4667), .Y(n6304) );
  AOI31X1 U9666 ( .A0(n6307), .A1(n6293), .A2(n6292), .B0(n6304), .Y(n6294) );
  NOR2BX1 U9667 ( .AN(n5936), .B(N3355), .Y(n6305) );
  NOR2X1 U9668 ( .A(n6150), .B(n6305), .Y(n6306) );
  AOI211X1 U9669 ( .A0(n6294), .A1(n6306), .B0(n6150), .C0(n6309), .Y(n6295)
         );
  NOR3BXL U9670 ( .AN(n6311), .B(n6310), .C(n6295), .Y(n6296) );
  NOR2X1 U9671 ( .A(n5950), .B(n5658), .Y(n6316) );
  AOI31X1 U9672 ( .A0(n6317), .A1(n6297), .A2(n6313), .B0(n6316), .Y(n6298) );
  OAI2BB1X1 U9673 ( .A0N(n6301), .A1N(n5922), .B0(N3358), .Y(n6300) );
  OAI211X1 U9674 ( .A0(n5921), .A1(n6301), .B0(n6300), .C0(n6299), .Y(n6303)
         );
  NAND3BX1 U9675 ( .AN(n6304), .B(n6303), .C(n6302), .Y(n6308) );
  AOI31X1 U9676 ( .A0(n6308), .A1(n6307), .A2(n6306), .B0(n6305), .Y(n6312) );
  AOI211X1 U9677 ( .A0(n6312), .A1(n6311), .B0(n6310), .C0(n6309), .Y(n6314)
         );
  OAI31XL U9678 ( .A0(n6316), .A1(n6315), .A2(n6314), .B0(n6313), .Y(N5603) );
  NAND2X1 U9679 ( .A(n5660), .B(n5946), .Y(n6326) );
  NAND2BX1 U9680 ( .AN(n5926), .B(n5664), .Y(n6321) );
  AO21X1 U9681 ( .A0(n5923), .A1(n6319), .B0(n5665), .Y(n6318) );
  NAND2BX1 U9682 ( .AN(n5664), .B(n5925), .Y(n6330) );
  OAI211X1 U9683 ( .A0(n6319), .A1(n5923), .B0(n6318), .C0(n6328), .Y(n6320)
         );
  NOR2X1 U9684 ( .A(n5931), .B(n5663), .Y(n6332) );
  NOR2BX1 U9685 ( .AN(n5662), .B(n5935), .Y(n6322) );
  NOR2BX1 U9686 ( .AN(n5936), .B(n5662), .Y(n6333) );
  NAND2X1 U9687 ( .A(N3360), .B(n5950), .Y(n6341) );
  NOR2X1 U9688 ( .A(n5950), .B(N3360), .Y(n6344) );
  OAI211X1 U9689 ( .A0(n5921), .A1(n6231), .B0(n6329), .C0(n6328), .Y(n6331)
         );
  NAND3BX1 U9690 ( .AN(n6332), .B(n6331), .C(n6330), .Y(n6336) );
  AOI31X1 U9691 ( .A0(n6336), .A1(n6335), .A2(n6334), .B0(n6333), .Y(n6340) );
  AOI211X1 U9692 ( .A0(n6340), .A1(n6339), .B0(n6338), .C0(n6337), .Y(n6342)
         );
endmodule

