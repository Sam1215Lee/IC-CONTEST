
module LCD_CTRL_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module LCD_CTRL_DW01_add_2 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [9:1] carry;

  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LCD_CTRL_DW01_add_1 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [9:1] carry;

  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module LCD_CTRL_DW01_add_0 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [9:1] carry;
  assign SUM[9] = carry[9];

  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  OAI2BB1X1 U1 ( .A0N(A[1]), .A1N(B[1]), .B0(n1), .Y(carry[2]) );
  OAI211X1 U2 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n1) );
endmodule


module LCD_CTRL ( clk, reset, IROM_Q, cmd, cmd_valid, IROM_EN, IROM_A, IRB_RW, 
        IRB_D, IRB_A, busy, done );
  input [7:0] IROM_Q;
  input [2:0] cmd;
  output [5:0] IROM_A;
  output [7:0] IRB_D;
  output [5:0] IRB_A;
  input clk, reset, cmd_valid;
  output IROM_EN, IRB_RW, busy, done;
  wire   N1656, N1657, N1658, N1659, N1661, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, \cnt[6] , \buff[0][7] , \buff[0][6] , \buff[0][5] ,
         \buff[0][4] , \buff[0][3] , \buff[0][2] , \buff[0][1] , \buff[0][0] ,
         \buff[1][7] , \buff[1][6] , \buff[1][5] , \buff[1][4] , \buff[1][3] ,
         \buff[1][2] , \buff[1][1] , \buff[1][0] , \buff[2][7] , \buff[2][6] ,
         \buff[2][5] , \buff[2][4] , \buff[2][3] , \buff[2][2] , \buff[2][1] ,
         \buff[2][0] , \buff[3][7] , \buff[3][6] , \buff[3][5] , \buff[3][4] ,
         \buff[3][3] , \buff[3][2] , \buff[3][1] , \buff[3][0] , \buff[4][7] ,
         \buff[4][6] , \buff[4][5] , \buff[4][4] , \buff[4][3] , \buff[4][2] ,
         \buff[4][1] , \buff[4][0] , \buff[5][7] , \buff[5][6] , \buff[5][5] ,
         \buff[5][4] , \buff[5][3] , \buff[5][2] , \buff[5][1] , \buff[5][0] ,
         \buff[6][7] , \buff[6][6] , \buff[6][5] , \buff[6][4] , \buff[6][3] ,
         \buff[6][2] , \buff[6][1] , \buff[6][0] , \buff[7][7] , \buff[7][6] ,
         \buff[7][5] , \buff[7][4] , \buff[7][3] , \buff[7][2] , \buff[7][1] ,
         \buff[7][0] , \buff[8][7] , \buff[8][6] , \buff[8][5] , \buff[8][4] ,
         \buff[8][3] , \buff[8][2] , \buff[8][1] , \buff[8][0] , \buff[9][7] ,
         \buff[9][6] , \buff[9][5] , \buff[9][4] , \buff[9][3] , \buff[9][2] ,
         \buff[9][1] , \buff[9][0] , \buff[10][7] , \buff[10][6] ,
         \buff[10][5] , \buff[10][4] , \buff[10][3] , \buff[10][2] ,
         \buff[10][1] , \buff[10][0] , \buff[11][7] , \buff[11][6] ,
         \buff[11][5] , \buff[11][4] , \buff[11][3] , \buff[11][2] ,
         \buff[11][1] , \buff[11][0] , \buff[12][7] , \buff[12][6] ,
         \buff[12][5] , \buff[12][4] , \buff[12][3] , \buff[12][2] ,
         \buff[12][1] , \buff[12][0] , \buff[13][7] , \buff[13][6] ,
         \buff[13][5] , \buff[13][4] , \buff[13][3] , \buff[13][2] ,
         \buff[13][1] , \buff[13][0] , \buff[14][7] , \buff[14][6] ,
         \buff[14][5] , \buff[14][4] , \buff[14][3] , \buff[14][2] ,
         \buff[14][1] , \buff[14][0] , \buff[15][7] , \buff[15][6] ,
         \buff[15][5] , \buff[15][4] , \buff[15][3] , \buff[15][2] ,
         \buff[15][1] , \buff[15][0] , \buff[16][7] , \buff[16][6] ,
         \buff[16][5] , \buff[16][4] , \buff[16][3] , \buff[16][2] ,
         \buff[16][1] , \buff[16][0] , \buff[17][7] , \buff[17][6] ,
         \buff[17][5] , \buff[17][4] , \buff[17][3] , \buff[17][2] ,
         \buff[17][1] , \buff[17][0] , \buff[18][7] , \buff[18][6] ,
         \buff[18][5] , \buff[18][4] , \buff[18][3] , \buff[18][2] ,
         \buff[18][1] , \buff[18][0] , \buff[19][7] , \buff[19][6] ,
         \buff[19][5] , \buff[19][4] , \buff[19][3] , \buff[19][2] ,
         \buff[19][1] , \buff[19][0] , \buff[20][7] , \buff[20][6] ,
         \buff[20][5] , \buff[20][4] , \buff[20][3] , \buff[20][2] ,
         \buff[20][1] , \buff[20][0] , \buff[21][7] , \buff[21][6] ,
         \buff[21][5] , \buff[21][4] , \buff[21][3] , \buff[21][2] ,
         \buff[21][1] , \buff[21][0] , \buff[22][7] , \buff[22][6] ,
         \buff[22][5] , \buff[22][4] , \buff[22][3] , \buff[22][2] ,
         \buff[22][1] , \buff[22][0] , \buff[23][7] , \buff[23][6] ,
         \buff[23][5] , \buff[23][4] , \buff[23][3] , \buff[23][2] ,
         \buff[23][1] , \buff[23][0] , \buff[24][7] , \buff[24][6] ,
         \buff[24][5] , \buff[24][4] , \buff[24][3] , \buff[24][2] ,
         \buff[24][1] , \buff[24][0] , \buff[25][7] , \buff[25][6] ,
         \buff[25][5] , \buff[25][4] , \buff[25][3] , \buff[25][2] ,
         \buff[25][1] , \buff[25][0] , \buff[26][7] , \buff[26][6] ,
         \buff[26][5] , \buff[26][4] , \buff[26][3] , \buff[26][2] ,
         \buff[26][1] , \buff[26][0] , \buff[27][7] , \buff[27][6] ,
         \buff[27][5] , \buff[27][4] , \buff[27][3] , \buff[27][2] ,
         \buff[27][1] , \buff[27][0] , \buff[28][7] , \buff[28][6] ,
         \buff[28][5] , \buff[28][4] , \buff[28][3] , \buff[28][2] ,
         \buff[28][1] , \buff[28][0] , \buff[29][7] , \buff[29][6] ,
         \buff[29][5] , \buff[29][4] , \buff[29][3] , \buff[29][2] ,
         \buff[29][1] , \buff[29][0] , \buff[30][7] , \buff[30][6] ,
         \buff[30][5] , \buff[30][4] , \buff[30][3] , \buff[30][2] ,
         \buff[30][1] , \buff[30][0] , \buff[31][7] , \buff[31][6] ,
         \buff[31][5] , \buff[31][4] , \buff[31][3] , \buff[31][2] ,
         \buff[31][1] , \buff[31][0] , \buff[32][7] , \buff[32][6] ,
         \buff[32][5] , \buff[32][4] , \buff[32][3] , \buff[32][2] ,
         \buff[32][1] , \buff[32][0] , \buff[33][7] , \buff[33][6] ,
         \buff[33][5] , \buff[33][4] , \buff[33][3] , \buff[33][2] ,
         \buff[33][1] , \buff[33][0] , \buff[34][7] , \buff[34][6] ,
         \buff[34][5] , \buff[34][4] , \buff[34][3] , \buff[34][2] ,
         \buff[34][1] , \buff[34][0] , \buff[35][7] , \buff[35][6] ,
         \buff[35][5] , \buff[35][4] , \buff[35][3] , \buff[35][2] ,
         \buff[35][1] , \buff[35][0] , \buff[36][7] , \buff[36][6] ,
         \buff[36][5] , \buff[36][4] , \buff[36][3] , \buff[36][2] ,
         \buff[36][1] , \buff[36][0] , \buff[37][7] , \buff[37][6] ,
         \buff[37][5] , \buff[37][4] , \buff[37][3] , \buff[37][2] ,
         \buff[37][1] , \buff[37][0] , \buff[38][7] , \buff[38][6] ,
         \buff[38][5] , \buff[38][4] , \buff[38][3] , \buff[38][2] ,
         \buff[38][1] , \buff[38][0] , \buff[39][7] , \buff[39][6] ,
         \buff[39][5] , \buff[39][4] , \buff[39][3] , \buff[39][2] ,
         \buff[39][1] , \buff[39][0] , \buff[40][7] , \buff[40][6] ,
         \buff[40][5] , \buff[40][4] , \buff[40][3] , \buff[40][2] ,
         \buff[40][1] , \buff[40][0] , \buff[41][7] , \buff[41][6] ,
         \buff[41][5] , \buff[41][4] , \buff[41][3] , \buff[41][2] ,
         \buff[41][1] , \buff[41][0] , \buff[42][7] , \buff[42][6] ,
         \buff[42][5] , \buff[42][4] , \buff[42][3] , \buff[42][2] ,
         \buff[42][1] , \buff[42][0] , \buff[43][7] , \buff[43][6] ,
         \buff[43][5] , \buff[43][4] , \buff[43][3] , \buff[43][2] ,
         \buff[43][1] , \buff[43][0] , \buff[44][7] , \buff[44][6] ,
         \buff[44][5] , \buff[44][4] , \buff[44][3] , \buff[44][2] ,
         \buff[44][1] , \buff[44][0] , \buff[45][7] , \buff[45][6] ,
         \buff[45][5] , \buff[45][4] , \buff[45][3] , \buff[45][2] ,
         \buff[45][1] , \buff[45][0] , \buff[46][7] , \buff[46][6] ,
         \buff[46][5] , \buff[46][4] , \buff[46][3] , \buff[46][2] ,
         \buff[46][1] , \buff[46][0] , \buff[47][7] , \buff[47][6] ,
         \buff[47][5] , \buff[47][4] , \buff[47][3] , \buff[47][2] ,
         \buff[47][1] , \buff[47][0] , \buff[48][7] , \buff[48][6] ,
         \buff[48][5] , \buff[48][4] , \buff[48][3] , \buff[48][2] ,
         \buff[48][1] , \buff[48][0] , \buff[49][7] , \buff[49][6] ,
         \buff[49][5] , \buff[49][4] , \buff[49][3] , \buff[49][2] ,
         \buff[49][1] , \buff[49][0] , \buff[50][7] , \buff[50][6] ,
         \buff[50][5] , \buff[50][4] , \buff[50][3] , \buff[50][2] ,
         \buff[50][1] , \buff[50][0] , \buff[51][7] , \buff[51][6] ,
         \buff[51][5] , \buff[51][4] , \buff[51][3] , \buff[51][2] ,
         \buff[51][1] , \buff[51][0] , \buff[52][7] , \buff[52][6] ,
         \buff[52][5] , \buff[52][4] , \buff[52][3] , \buff[52][2] ,
         \buff[52][1] , \buff[52][0] , \buff[53][7] , \buff[53][6] ,
         \buff[53][5] , \buff[53][4] , \buff[53][3] , \buff[53][2] ,
         \buff[53][1] , \buff[53][0] , \buff[54][7] , \buff[54][6] ,
         \buff[54][5] , \buff[54][4] , \buff[54][3] , \buff[54][2] ,
         \buff[54][1] , \buff[54][0] , \buff[55][7] , \buff[55][6] ,
         \buff[55][5] , \buff[55][4] , \buff[55][3] , \buff[55][2] ,
         \buff[55][1] , \buff[55][0] , \buff[56][7] , \buff[56][6] ,
         \buff[56][5] , \buff[56][4] , \buff[56][3] , \buff[56][2] ,
         \buff[56][1] , \buff[56][0] , \buff[57][7] , \buff[57][6] ,
         \buff[57][5] , \buff[57][4] , \buff[57][3] , \buff[57][2] ,
         \buff[57][1] , \buff[57][0] , \buff[58][7] , \buff[58][6] ,
         \buff[58][5] , \buff[58][4] , \buff[58][3] , \buff[58][2] ,
         \buff[58][1] , \buff[58][0] , \buff[59][7] , \buff[59][6] ,
         \buff[59][5] , \buff[59][4] , \buff[59][3] , \buff[59][2] ,
         \buff[59][1] , \buff[59][0] , \buff[60][7] , \buff[60][6] ,
         \buff[60][5] , \buff[60][4] , \buff[60][3] , \buff[60][2] ,
         \buff[60][1] , \buff[60][0] , \buff[61][7] , \buff[61][6] ,
         \buff[61][5] , \buff[61][4] , \buff[61][3] , \buff[61][2] ,
         \buff[61][1] , \buff[61][0] , \buff[62][7] , \buff[62][6] ,
         \buff[62][5] , \buff[62][4] , \buff[62][3] , \buff[62][2] ,
         \buff[62][1] , \buff[62][0] , \buff[63][7] , \buff[63][6] ,
         \buff[63][5] , \buff[63][4] , \buff[63][3] , \buff[63][2] ,
         \buff[63][1] , \buff[63][0] , N1677, N1743, N1744, N1745, N1746,
         N1747, N1748, N1749, N7371, N7372, N7373, N7374, N7375, N7376, N7377,
         N7378, N7380, N7381, N7382, N7383, N7384, N7385, N7386, N7387, N7388,
         N7391, N7392, N7393, N7395, n91, n92, n94, n96, n98, n99, n100, n101,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n148, n149,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n238, n240, n241, n243, n244, n245, n246,
         n250, n251, n252, n253, n257, n258, n259, n260, n264, n265, n266,
         n267, n271, n272, n273, n274, n278, n279, n280, n281, n285, n286,
         n287, n288, n292, n293, n296, n298, n299, n301, n302, n304, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n317, n318,
         n320, n321, n322, n323, n325, n326, n328, n329, n330, n331, n333,
         n334, n336, n337, n338, n339, n341, n342, n344, n345, n346, n347,
         n349, n350, n351, n352, n353, n354, n355, n357, n358, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n370, n371, n373, n374,
         n375, n376, n377, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n667, n668, n669,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n709, n710, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n748, n749, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n787, n788, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n826, n827, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n865, n866,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n904, n905, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n985, n988, n989, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1029, n1030, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1068, n1069, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1107, n1108, n1110,
         n1111, n1112, n1113, n1114, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1146, n1147, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1185, n1186, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1224, n1225, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1303, n1304, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1344, n1345, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1383,
         n1384, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1459, n1461, n1463, n1464, n1466, n1467, n1468,
         n1469, n1470, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1502, n1503, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1541, n1542,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1619, n1620, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1659, n1660, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1698,
         n1699, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1737, n1738, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1817, n1818, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1856, n1857,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1972, n1973, n1974, n1975, n1976, n1977, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2015, n2016, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2054,
         n2055, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2093, n2094, n2096, n2097,
         n2098, n2099, n2100, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2132, n2133, n2134, n2136, n2137, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2175, n2176, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2254, n2255, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2298,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2335, n2336, n2338, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2375, n2376, n2378, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2453, n2454, n2455, n2456,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2494, n2495, n2497, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2535, n2536, n2538, n2539, n2540, n2541, n2544,
         n2546, n2547, n2549, n2550, n2551, n2552, n2555, n2557, n2558, n2559,
         n2560, n2562, n2563, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, N7429, N7428, N7427, N7426, N7425, N7424, N7423,
         N7422, N7421, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8393, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825;
  wire   [1:0] next;
  wire   [9:2] avg_reg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign done = 1'b1;

  OAI221X2 U214 ( .A0(n9613), .A1(n9796), .B0(n9608), .B1(n9789), .C0(n9663), 
        .Y(n238) );
  OAI211X2 U2997 ( .A0(IRB_RW), .A1(n91), .B0(n2567), .C0(n2568), .Y(n2566) );
  LCD_CTRL_DW01_inc_0 r1252 ( .A({\cnt[6] , N1661, n8393, N1659, N1658, N1657, 
        n9317}), .SUM({N1749, N1748, N1747, N1746, N1745, N1744, N1743}) );
  LCD_CTRL_DW01_add_2 add_2_root_add_0_root_add_170_3 ( .A({1'b0, 1'b0, N7380, 
        N7381, N7382, N7383, N7384, N7385, N7386, N7387}), .B({1'b0, 1'b0, 
        n7231, n7230, n7229, n7228, n7234, n7227, n8420, n8419}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N7429, N7428, N7427, N7426, N7425, 
        N7424, N7423, N7422, N7421}) );
  LCD_CTRL_DW01_add_1 add_1_root_add_0_root_add_170_3 ( .A({1'b0, 1'b0, N7395, 
        n7235, N7393, N7392, N7391, n7233, n8418, N7388}), .B({1'b0, 1'b0, 
        n8445, n8444, n8443, n8442, n8435, n8434, n8437, n8436}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__1, n9825, n9824, n9823, n9822, n9821, 
        n9820, n9819, n9818, n9817}) );
  LCD_CTRL_DW01_add_0 add_0_root_add_0_root_add_170_3 ( .A({1'b0, N7429, N7428, 
        N7427, N7426, N7425, N7424, N7423, N7422, N7421}), .B({1'b0, n9825, 
        n9824, n9823, n9822, n9821, n9820, n9819, n9818, n9817}), .CI(1'b0), 
        .SUM({avg_reg, SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3}) );
  DFFQX1 \buff_reg[63][7]  ( .D(n8336), .CK(clk), .Q(\buff[63][7] ) );
  DFFQX1 \buff_reg[63][6]  ( .D(n8361), .CK(clk), .Q(\buff[63][6] ) );
  DFFQX1 \buff_reg[63][5]  ( .D(n7267), .CK(clk), .Q(\buff[63][5] ) );
  DFFQX1 \buff_reg[63][4]  ( .D(n7266), .CK(clk), .Q(\buff[63][4] ) );
  DFFQX1 \buff_reg[63][3]  ( .D(n7261), .CK(clk), .Q(\buff[63][3] ) );
  DFFQX1 \buff_reg[63][2]  ( .D(n7258), .CK(clk), .Q(\buff[63][2] ) );
  DFFQX1 \buff_reg[63][1]  ( .D(n7255), .CK(clk), .Q(\buff[63][1] ) );
  DFFQX1 \buff_reg[63][0]  ( .D(n7252), .CK(clk), .Q(\buff[63][0] ) );
  DFFQX1 \buff_reg[61][7]  ( .D(n2617), .CK(clk), .Q(\buff[61][7] ) );
  DFFQX1 \buff_reg[61][6]  ( .D(n2616), .CK(clk), .Q(\buff[61][6] ) );
  DFFQX1 \buff_reg[61][5]  ( .D(n2615), .CK(clk), .Q(\buff[61][5] ) );
  DFFQX1 \buff_reg[61][4]  ( .D(n7312), .CK(clk), .Q(\buff[61][4] ) );
  DFFQX1 \buff_reg[61][3]  ( .D(n7309), .CK(clk), .Q(\buff[61][3] ) );
  DFFQX1 \buff_reg[61][2]  ( .D(n7306), .CK(clk), .Q(\buff[61][2] ) );
  DFFQX1 \buff_reg[61][1]  ( .D(n7303), .CK(clk), .Q(\buff[61][1] ) );
  DFFQX1 \buff_reg[61][0]  ( .D(n7300), .CK(clk), .Q(\buff[61][0] ) );
  DFFQX1 \buff_reg[59][7]  ( .D(n7297), .CK(clk), .Q(\buff[59][7] ) );
  DFFQX1 \buff_reg[59][6]  ( .D(n2632), .CK(clk), .Q(\buff[59][6] ) );
  DFFQX1 \buff_reg[59][5]  ( .D(n7363), .CK(clk), .Q(\buff[59][5] ) );
  DFFQX1 \buff_reg[59][4]  ( .D(n7362), .CK(clk), .Q(\buff[59][4] ) );
  DFFQX1 \buff_reg[59][3]  ( .D(n7357), .CK(clk), .Q(\buff[59][3] ) );
  DFFQX1 \buff_reg[59][2]  ( .D(n7354), .CK(clk), .Q(\buff[59][2] ) );
  DFFQX1 \buff_reg[59][1]  ( .D(n7351), .CK(clk), .Q(\buff[59][1] ) );
  DFFQX1 \buff_reg[59][0]  ( .D(n7348), .CK(clk), .Q(\buff[59][0] ) );
  DFFQX1 \buff_reg[57][7]  ( .D(n2649), .CK(clk), .Q(\buff[57][7] ) );
  DFFQX1 \buff_reg[57][6]  ( .D(n2648), .CK(clk), .Q(\buff[57][6] ) );
  DFFQX1 \buff_reg[57][5]  ( .D(n2647), .CK(clk), .Q(\buff[57][5] ) );
  DFFQX1 \buff_reg[57][4]  ( .D(n7406), .CK(clk), .Q(\buff[57][4] ) );
  DFFQX1 \buff_reg[57][3]  ( .D(n7403), .CK(clk), .Q(\buff[57][3] ) );
  DFFQX1 \buff_reg[57][2]  ( .D(n7400), .CK(clk), .Q(\buff[57][2] ) );
  DFFQX1 \buff_reg[57][1]  ( .D(n7397), .CK(clk), .Q(\buff[57][1] ) );
  DFFQX1 \buff_reg[57][0]  ( .D(n7394), .CK(clk), .Q(\buff[57][0] ) );
  DFFQX1 \buff_reg[60][7]  ( .D(n2625), .CK(clk), .Q(\buff[60][7] ) );
  DFFQX1 \buff_reg[60][6]  ( .D(n2624), .CK(clk), .Q(\buff[60][6] ) );
  DFFQX1 \buff_reg[60][5]  ( .D(n2623), .CK(clk), .Q(\buff[60][5] ) );
  DFFQX1 \buff_reg[60][4]  ( .D(n7336), .CK(clk), .Q(\buff[60][4] ) );
  DFFQX1 \buff_reg[60][3]  ( .D(n7333), .CK(clk), .Q(\buff[60][3] ) );
  DFFQX1 \buff_reg[60][2]  ( .D(n7330), .CK(clk), .Q(\buff[60][2] ) );
  DFFQX1 \buff_reg[60][1]  ( .D(n7327), .CK(clk), .Q(\buff[60][1] ) );
  DFFQX1 \buff_reg[60][0]  ( .D(n7324), .CK(clk), .Q(\buff[60][0] ) );
  DFFQX1 \buff_reg[62][7]  ( .D(n2609), .CK(clk), .Q(\buff[62][7] ) );
  DFFQX1 \buff_reg[62][6]  ( .D(n2608), .CK(clk), .Q(\buff[62][6] ) );
  DFFQX1 \buff_reg[62][5]  ( .D(n2607), .CK(clk), .Q(\buff[62][5] ) );
  DFFQX1 \buff_reg[62][4]  ( .D(n7288), .CK(clk), .Q(\buff[62][4] ) );
  DFFQX1 \buff_reg[62][3]  ( .D(n7285), .CK(clk), .Q(\buff[62][3] ) );
  DFFQX1 \buff_reg[62][2]  ( .D(n7282), .CK(clk), .Q(\buff[62][2] ) );
  DFFQX1 \buff_reg[62][1]  ( .D(n7279), .CK(clk), .Q(\buff[62][1] ) );
  DFFQX1 \buff_reg[62][0]  ( .D(n7276), .CK(clk), .Q(\buff[62][0] ) );
  DFFQX1 \buff_reg[56][7]  ( .D(n2657), .CK(clk), .Q(\buff[56][7] ) );
  DFFQX1 \buff_reg[56][6]  ( .D(n2656), .CK(clk), .Q(\buff[56][6] ) );
  DFFQX1 \buff_reg[56][5]  ( .D(n2655), .CK(clk), .Q(\buff[56][5] ) );
  DFFQX1 \buff_reg[56][4]  ( .D(n7430), .CK(clk), .Q(\buff[56][4] ) );
  DFFQX1 \buff_reg[56][3]  ( .D(n7427), .CK(clk), .Q(\buff[56][3] ) );
  DFFQX1 \buff_reg[56][2]  ( .D(n7424), .CK(clk), .Q(\buff[56][2] ) );
  DFFQX1 \buff_reg[56][1]  ( .D(n7421), .CK(clk), .Q(\buff[56][1] ) );
  DFFQX1 \buff_reg[56][0]  ( .D(n7418), .CK(clk), .Q(\buff[56][0] ) );
  DFFQX1 \buff_reg[58][7]  ( .D(n2641), .CK(clk), .Q(\buff[58][7] ) );
  DFFQX1 \buff_reg[58][6]  ( .D(n2640), .CK(clk), .Q(\buff[58][6] ) );
  DFFQX1 \buff_reg[58][5]  ( .D(n2639), .CK(clk), .Q(\buff[58][5] ) );
  DFFQX1 \buff_reg[58][4]  ( .D(n7382), .CK(clk), .Q(\buff[58][4] ) );
  DFFQX1 \buff_reg[58][3]  ( .D(n7379), .CK(clk), .Q(\buff[58][3] ) );
  DFFQX1 \buff_reg[58][2]  ( .D(n7376), .CK(clk), .Q(\buff[58][2] ) );
  DFFQX1 \buff_reg[58][1]  ( .D(n7373), .CK(clk), .Q(\buff[58][1] ) );
  DFFQX1 \buff_reg[58][0]  ( .D(n7370), .CK(clk), .Q(\buff[58][0] ) );
  DFFQX1 \buff_reg[28][7]  ( .D(n2881), .CK(clk), .Q(\buff[28][7] ) );
  DFFQX1 \buff_reg[28][6]  ( .D(n2880), .CK(clk), .Q(\buff[28][6] ) );
  DFFQX1 \buff_reg[28][5]  ( .D(n7880), .CK(clk), .Q(\buff[28][5] ) );
  DFFQX1 \buff_reg[28][4]  ( .D(n7878), .CK(clk), .Q(\buff[28][4] ) );
  DFFQX1 \buff_reg[28][3]  ( .D(n7876), .CK(clk), .Q(\buff[28][3] ) );
  DFFQX1 \buff_reg[28][2]  ( .D(n7874), .CK(clk), .Q(\buff[28][2] ) );
  DFFQX1 \buff_reg[28][1]  ( .D(n7872), .CK(clk), .Q(\buff[28][1] ) );
  DFFQX1 \buff_reg[28][0]  ( .D(n7870), .CK(clk), .Q(\buff[28][0] ) );
  DFFQX1 \buff_reg[30][7]  ( .D(n2865), .CK(clk), .Q(\buff[30][7] ) );
  DFFQX1 \buff_reg[30][6]  ( .D(n2864), .CK(clk), .Q(\buff[30][6] ) );
  DFFQX1 \buff_reg[30][5]  ( .D(n7848), .CK(clk), .Q(\buff[30][5] ) );
  DFFQX1 \buff_reg[30][4]  ( .D(n7846), .CK(clk), .Q(\buff[30][4] ) );
  DFFQX1 \buff_reg[30][3]  ( .D(n7844), .CK(clk), .Q(\buff[30][3] ) );
  DFFQX1 \buff_reg[30][2]  ( .D(n7842), .CK(clk), .Q(\buff[30][2] ) );
  DFFQX1 \buff_reg[30][1]  ( .D(n7840), .CK(clk), .Q(\buff[30][1] ) );
  DFFQX1 \buff_reg[30][0]  ( .D(n7838), .CK(clk), .Q(\buff[30][0] ) );
  DFFQX1 \buff_reg[24][7]  ( .D(n2913), .CK(clk), .Q(\buff[24][7] ) );
  DFFQX1 \buff_reg[24][6]  ( .D(n2912), .CK(clk), .Q(\buff[24][6] ) );
  DFFQX1 \buff_reg[24][5]  ( .D(n7944), .CK(clk), .Q(\buff[24][5] ) );
  DFFQX1 \buff_reg[24][4]  ( .D(n7942), .CK(clk), .Q(\buff[24][4] ) );
  DFFQX1 \buff_reg[24][3]  ( .D(n7940), .CK(clk), .Q(\buff[24][3] ) );
  DFFQX1 \buff_reg[24][2]  ( .D(n7938), .CK(clk), .Q(\buff[24][2] ) );
  DFFQX1 \buff_reg[24][1]  ( .D(n7936), .CK(clk), .Q(\buff[24][1] ) );
  DFFQX1 \buff_reg[24][0]  ( .D(n7934), .CK(clk), .Q(\buff[24][0] ) );
  DFFQX1 \buff_reg[26][7]  ( .D(n2897), .CK(clk), .Q(\buff[26][7] ) );
  DFFQX1 \buff_reg[26][6]  ( .D(n2896), .CK(clk), .Q(\buff[26][6] ) );
  DFFQX1 \buff_reg[26][5]  ( .D(n2895), .CK(clk), .Q(\buff[26][5] ) );
  DFFQX1 \buff_reg[26][4]  ( .D(n2894), .CK(clk), .Q(\buff[26][4] ) );
  DFFQX1 \buff_reg[26][3]  ( .D(n2893), .CK(clk), .Q(\buff[26][3] ) );
  DFFQX1 \buff_reg[26][2]  ( .D(n2892), .CK(clk), .Q(\buff[26][2] ) );
  DFFQX1 \buff_reg[26][1]  ( .D(n2891), .CK(clk), .Q(\buff[26][1] ) );
  DFFQX1 \buff_reg[26][0]  ( .D(n7902), .CK(clk), .Q(\buff[26][0] ) );
  DFFQX1 \buff_reg[4][7]  ( .D(n3073), .CK(clk), .Q(\buff[4][7] ) );
  DFFQX1 \buff_reg[4][6]  ( .D(n3072), .CK(clk), .Q(\buff[4][6] ) );
  DFFQX1 \buff_reg[4][5]  ( .D(n8268), .CK(clk), .Q(\buff[4][5] ) );
  DFFQX1 \buff_reg[4][4]  ( .D(n8266), .CK(clk), .Q(\buff[4][4] ) );
  DFFQX1 \buff_reg[4][3]  ( .D(n3069), .CK(clk), .Q(\buff[4][3] ) );
  DFFQX1 \buff_reg[4][2]  ( .D(n8261), .CK(clk), .Q(\buff[4][2] ) );
  DFFQX1 \buff_reg[4][1]  ( .D(n8259), .CK(clk), .Q(\buff[4][1] ) );
  DFFQX1 \buff_reg[4][0]  ( .D(n8257), .CK(clk), .Q(\buff[4][0] ) );
  DFFQX1 \buff_reg[12][7]  ( .D(n3009), .CK(clk), .Q(\buff[12][7] ) );
  DFFQX1 \buff_reg[12][6]  ( .D(n3008), .CK(clk), .Q(\buff[12][6] ) );
  DFFQX1 \buff_reg[12][5]  ( .D(n8137), .CK(clk), .Q(\buff[12][5] ) );
  DFFQX1 \buff_reg[12][4]  ( .D(n8135), .CK(clk), .Q(\buff[12][4] ) );
  DFFQX1 \buff_reg[12][3]  ( .D(n8133), .CK(clk), .Q(\buff[12][3] ) );
  DFFQX1 \buff_reg[12][2]  ( .D(n8131), .CK(clk), .Q(\buff[12][2] ) );
  DFFQX1 \buff_reg[12][1]  ( .D(n8129), .CK(clk), .Q(\buff[12][1] ) );
  DFFQX1 \buff_reg[12][0]  ( .D(n8127), .CK(clk), .Q(\buff[12][0] ) );
  DFFQX1 \buff_reg[20][7]  ( .D(n2945), .CK(clk), .Q(\buff[20][7] ) );
  DFFQX1 \buff_reg[20][6]  ( .D(n2944), .CK(clk), .Q(\buff[20][6] ) );
  DFFQX1 \buff_reg[20][5]  ( .D(n8008), .CK(clk), .Q(\buff[20][5] ) );
  DFFQX1 \buff_reg[20][4]  ( .D(n8006), .CK(clk), .Q(\buff[20][4] ) );
  DFFQX1 \buff_reg[20][3]  ( .D(n8004), .CK(clk), .Q(\buff[20][3] ) );
  DFFQX1 \buff_reg[20][2]  ( .D(n8002), .CK(clk), .Q(\buff[20][2] ) );
  DFFQX1 \buff_reg[20][1]  ( .D(n8000), .CK(clk), .Q(\buff[20][1] ) );
  DFFQX1 \buff_reg[20][0]  ( .D(n7998), .CK(clk), .Q(\buff[20][0] ) );
  DFFQX1 \buff_reg[36][7]  ( .D(n7996), .CK(clk), .Q(\buff[36][7] ) );
  DFFQX1 \buff_reg[36][6]  ( .D(n7994), .CK(clk), .Q(\buff[36][6] ) );
  DFFQX1 \buff_reg[36][5]  ( .D(n7751), .CK(clk), .Q(\buff[36][5] ) );
  DFFQX1 \buff_reg[36][4]  ( .D(n7749), .CK(clk), .Q(\buff[36][4] ) );
  DFFQX1 \buff_reg[36][3]  ( .D(n7747), .CK(clk), .Q(\buff[36][3] ) );
  DFFQX1 \buff_reg[36][2]  ( .D(n7745), .CK(clk), .Q(\buff[36][2] ) );
  DFFQX1 \buff_reg[36][1]  ( .D(n7743), .CK(clk), .Q(\buff[36][1] ) );
  DFFQX1 \buff_reg[36][0]  ( .D(n7741), .CK(clk), .Q(\buff[36][0] ) );
  DFFQX1 \buff_reg[44][7]  ( .D(n2753), .CK(clk), .Q(\buff[44][7] ) );
  DFFQX1 \buff_reg[44][6]  ( .D(n2752), .CK(clk), .Q(\buff[44][6] ) );
  DFFQX1 \buff_reg[44][5]  ( .D(n7623), .CK(clk), .Q(\buff[44][5] ) );
  DFFQX1 \buff_reg[44][4]  ( .D(n7621), .CK(clk), .Q(\buff[44][4] ) );
  DFFQX1 \buff_reg[44][3]  ( .D(n7619), .CK(clk), .Q(\buff[44][3] ) );
  DFFQX1 \buff_reg[44][2]  ( .D(n7617), .CK(clk), .Q(\buff[44][2] ) );
  DFFQX1 \buff_reg[44][1]  ( .D(n7615), .CK(clk), .Q(\buff[44][1] ) );
  DFFQX1 \buff_reg[44][0]  ( .D(n7613), .CK(clk), .Q(\buff[44][0] ) );
  DFFQX1 \buff_reg[52][7]  ( .D(n7611), .CK(clk), .Q(\buff[52][7] ) );
  DFFQX1 \buff_reg[52][6]  ( .D(n7609), .CK(clk), .Q(\buff[52][6] ) );
  DFFQX1 \buff_reg[52][5]  ( .D(n7497), .CK(clk), .Q(\buff[52][5] ) );
  DFFQX1 \buff_reg[52][4]  ( .D(n7495), .CK(clk), .Q(\buff[52][4] ) );
  DFFQX1 \buff_reg[52][3]  ( .D(n7493), .CK(clk), .Q(\buff[52][3] ) );
  DFFQX1 \buff_reg[52][2]  ( .D(n2684), .CK(clk), .Q(\buff[52][2] ) );
  DFFQX1 \buff_reg[52][1]  ( .D(n2683), .CK(clk), .Q(\buff[52][1] ) );
  DFFQX1 \buff_reg[52][0]  ( .D(n7487), .CK(clk), .Q(\buff[52][0] ) );
  DFFQX1 \buff_reg[6][7]  ( .D(n3057), .CK(clk), .Q(\buff[6][7] ) );
  DFFQX1 \buff_reg[6][6]  ( .D(n3056), .CK(clk), .Q(\buff[6][6] ) );
  DFFQX1 \buff_reg[6][5]  ( .D(n3055), .CK(clk), .Q(\buff[6][5] ) );
  DFFQX1 \buff_reg[6][4]  ( .D(n3054), .CK(clk), .Q(\buff[6][4] ) );
  DFFQX1 \buff_reg[6][3]  ( .D(n3053), .CK(clk), .Q(\buff[6][3] ) );
  DFFQX1 \buff_reg[6][2]  ( .D(n3052), .CK(clk), .Q(\buff[6][2] ) );
  DFFQX1 \buff_reg[6][1]  ( .D(n3051), .CK(clk), .Q(\buff[6][1] ) );
  DFFQX1 \buff_reg[6][0]  ( .D(n3050), .CK(clk), .Q(\buff[6][0] ) );
  DFFQX1 \buff_reg[14][7]  ( .D(n8223), .CK(clk), .Q(\buff[14][7] ) );
  DFFQX1 \buff_reg[14][6]  ( .D(n2992), .CK(clk), .Q(\buff[14][6] ) );
  DFFQX1 \buff_reg[14][5]  ( .D(n8105), .CK(clk), .Q(\buff[14][5] ) );
  DFFQX1 \buff_reg[14][4]  ( .D(n8102), .CK(clk), .Q(\buff[14][4] ) );
  DFFQX1 \buff_reg[14][3]  ( .D(n8100), .CK(clk), .Q(\buff[14][3] ) );
  DFFQX1 \buff_reg[14][2]  ( .D(n8098), .CK(clk), .Q(\buff[14][2] ) );
  DFFQX1 \buff_reg[14][1]  ( .D(n8096), .CK(clk), .Q(\buff[14][1] ) );
  DFFQX1 \buff_reg[14][0]  ( .D(n8094), .CK(clk), .Q(\buff[14][0] ) );
  DFFQX1 \buff_reg[22][7]  ( .D(n2929), .CK(clk), .Q(\buff[22][7] ) );
  DFFQX1 \buff_reg[22][6]  ( .D(n2928), .CK(clk), .Q(\buff[22][6] ) );
  DFFQX1 \buff_reg[22][5]  ( .D(n7976), .CK(clk), .Q(\buff[22][5] ) );
  DFFQX1 \buff_reg[22][4]  ( .D(n7974), .CK(clk), .Q(\buff[22][4] ) );
  DFFQX1 \buff_reg[22][3]  ( .D(n7972), .CK(clk), .Q(\buff[22][3] ) );
  DFFQX1 \buff_reg[22][2]  ( .D(n7970), .CK(clk), .Q(\buff[22][2] ) );
  DFFQX1 \buff_reg[22][1]  ( .D(n7968), .CK(clk), .Q(\buff[22][1] ) );
  DFFQX1 \buff_reg[22][0]  ( .D(n7966), .CK(clk), .Q(\buff[22][0] ) );
  DFFQX1 \buff_reg[38][7]  ( .D(n7964), .CK(clk), .Q(\buff[38][7] ) );
  DFFQX1 \buff_reg[38][6]  ( .D(n7962), .CK(clk), .Q(\buff[38][6] ) );
  DFFQX1 \buff_reg[38][5]  ( .D(n7719), .CK(clk), .Q(\buff[38][5] ) );
  DFFQX1 \buff_reg[38][4]  ( .D(n7717), .CK(clk), .Q(\buff[38][4] ) );
  DFFQX1 \buff_reg[38][3]  ( .D(n7715), .CK(clk), .Q(\buff[38][3] ) );
  DFFQX1 \buff_reg[38][2]  ( .D(n7713), .CK(clk), .Q(\buff[38][2] ) );
  DFFQX1 \buff_reg[38][1]  ( .D(n7711), .CK(clk), .Q(\buff[38][1] ) );
  DFFQX1 \buff_reg[38][0]  ( .D(n7709), .CK(clk), .Q(\buff[38][0] ) );
  DFFQX1 \buff_reg[46][7]  ( .D(n2737), .CK(clk), .Q(\buff[46][7] ) );
  DFFQX1 \buff_reg[46][6]  ( .D(n2736), .CK(clk), .Q(\buff[46][6] ) );
  DFFQX1 \buff_reg[46][5]  ( .D(n7591), .CK(clk), .Q(\buff[46][5] ) );
  DFFQX1 \buff_reg[46][4]  ( .D(n7589), .CK(clk), .Q(\buff[46][4] ) );
  DFFQX1 \buff_reg[46][3]  ( .D(n7587), .CK(clk), .Q(\buff[46][3] ) );
  DFFQX1 \buff_reg[46][2]  ( .D(n7585), .CK(clk), .Q(\buff[46][2] ) );
  DFFQX1 \buff_reg[46][1]  ( .D(n7583), .CK(clk), .Q(\buff[46][1] ) );
  DFFQX1 \buff_reg[46][0]  ( .D(n7581), .CK(clk), .Q(\buff[46][0] ) );
  DFFQX1 \buff_reg[54][7]  ( .D(n7579), .CK(clk), .Q(\buff[54][7] ) );
  DFFQX1 \buff_reg[54][6]  ( .D(n7577), .CK(clk), .Q(\buff[54][6] ) );
  DFFQX1 \buff_reg[54][5]  ( .D(n7464), .CK(clk), .Q(\buff[54][5] ) );
  DFFQX1 \buff_reg[54][4]  ( .D(n7462), .CK(clk), .Q(\buff[54][4] ) );
  DFFQX1 \buff_reg[54][3]  ( .D(n7460), .CK(clk), .Q(\buff[54][3] ) );
  DFFQX1 \buff_reg[54][2]  ( .D(n7458), .CK(clk), .Q(\buff[54][2] ) );
  DFFQX1 \buff_reg[54][1]  ( .D(n7456), .CK(clk), .Q(\buff[54][1] ) );
  DFFQX1 \buff_reg[54][0]  ( .D(n7454), .CK(clk), .Q(\buff[54][0] ) );
  DFFQX1 \buff_reg[0][7]  ( .D(n3105), .CK(clk), .Q(\buff[0][7] ) );
  DFFQX1 \buff_reg[0][6]  ( .D(n3104), .CK(clk), .Q(\buff[0][6] ) );
  DFFQX1 \buff_reg[0][5]  ( .D(n8334), .CK(clk), .Q(\buff[0][5] ) );
  DFFQX1 \buff_reg[0][4]  ( .D(n8332), .CK(clk), .Q(\buff[0][4] ) );
  DFFQX1 \buff_reg[0][3]  ( .D(n3101), .CK(clk), .Q(\buff[0][3] ) );
  DFFQX1 \buff_reg[0][2]  ( .D(n8327), .CK(clk), .Q(\buff[0][2] ) );
  DFFQX1 \buff_reg[0][1]  ( .D(n8325), .CK(clk), .Q(\buff[0][1] ) );
  DFFQX1 \buff_reg[0][0]  ( .D(n8323), .CK(clk), .Q(\buff[0][0] ) );
  DFFQX1 \buff_reg[8][7]  ( .D(n8321), .CK(clk), .Q(\buff[8][7] ) );
  DFFQX1 \buff_reg[8][6]  ( .D(n3040), .CK(clk), .Q(\buff[8][6] ) );
  DFFQX1 \buff_reg[8][5]  ( .D(n8202), .CK(clk), .Q(\buff[8][5] ) );
  DFFQX1 \buff_reg[8][4]  ( .D(n8200), .CK(clk), .Q(\buff[8][4] ) );
  DFFQX1 \buff_reg[8][3]  ( .D(n8198), .CK(clk), .Q(\buff[8][3] ) );
  DFFQX1 \buff_reg[8][2]  ( .D(n8196), .CK(clk), .Q(\buff[8][2] ) );
  DFFQX1 \buff_reg[8][1]  ( .D(n8194), .CK(clk), .Q(\buff[8][1] ) );
  DFFQX1 \buff_reg[8][0]  ( .D(n8192), .CK(clk), .Q(\buff[8][0] ) );
  DFFQX1 \buff_reg[16][7]  ( .D(n8190), .CK(clk), .Q(\buff[16][7] ) );
  DFFQX1 \buff_reg[16][6]  ( .D(n2976), .CK(clk), .Q(\buff[16][6] ) );
  DFFQX1 \buff_reg[16][5]  ( .D(n8072), .CK(clk), .Q(\buff[16][5] ) );
  DFFQX1 \buff_reg[16][4]  ( .D(n8070), .CK(clk), .Q(\buff[16][4] ) );
  DFFQX1 \buff_reg[16][3]  ( .D(n8068), .CK(clk), .Q(\buff[16][3] ) );
  DFFQX1 \buff_reg[16][2]  ( .D(n8066), .CK(clk), .Q(\buff[16][2] ) );
  DFFQX1 \buff_reg[16][1]  ( .D(n8064), .CK(clk), .Q(\buff[16][1] ) );
  DFFQX1 \buff_reg[16][0]  ( .D(n8062), .CK(clk), .Q(\buff[16][0] ) );
  DFFQX1 \buff_reg[32][7]  ( .D(n8060), .CK(clk), .Q(\buff[32][7] ) );
  DFFQX1 \buff_reg[32][6]  ( .D(n8058), .CK(clk), .Q(\buff[32][6] ) );
  DFFQX1 \buff_reg[32][5]  ( .D(n7816), .CK(clk), .Q(\buff[32][5] ) );
  DFFQX1 \buff_reg[32][4]  ( .D(n7814), .CK(clk), .Q(\buff[32][4] ) );
  DFFQX1 \buff_reg[32][3]  ( .D(n7812), .CK(clk), .Q(\buff[32][3] ) );
  DFFQX1 \buff_reg[32][2]  ( .D(n7810), .CK(clk), .Q(\buff[32][2] ) );
  DFFQX1 \buff_reg[32][1]  ( .D(n2843), .CK(clk), .Q(\buff[32][1] ) );
  DFFQX1 \buff_reg[32][0]  ( .D(n7805), .CK(clk), .Q(\buff[32][0] ) );
  DFFQX1 \buff_reg[40][7]  ( .D(n2785), .CK(clk), .Q(\buff[40][7] ) );
  DFFQX1 \buff_reg[40][6]  ( .D(n2784), .CK(clk), .Q(\buff[40][6] ) );
  DFFQX1 \buff_reg[40][5]  ( .D(n7687), .CK(clk), .Q(\buff[40][5] ) );
  DFFQX1 \buff_reg[40][4]  ( .D(n7685), .CK(clk), .Q(\buff[40][4] ) );
  DFFQX1 \buff_reg[40][3]  ( .D(n7683), .CK(clk), .Q(\buff[40][3] ) );
  DFFQX1 \buff_reg[40][2]  ( .D(n7681), .CK(clk), .Q(\buff[40][2] ) );
  DFFQX1 \buff_reg[40][1]  ( .D(n7679), .CK(clk), .Q(\buff[40][1] ) );
  DFFQX1 \buff_reg[40][0]  ( .D(n7677), .CK(clk), .Q(\buff[40][0] ) );
  DFFQX1 \buff_reg[48][7]  ( .D(n7675), .CK(clk), .Q(\buff[48][7] ) );
  DFFQX1 \buff_reg[48][6]  ( .D(n7673), .CK(clk), .Q(\buff[48][6] ) );
  DFFQX1 \buff_reg[48][5]  ( .D(n7559), .CK(clk), .Q(\buff[48][5] ) );
  DFFQX1 \buff_reg[48][4]  ( .D(n7557), .CK(clk), .Q(\buff[48][4] ) );
  DFFQX1 \buff_reg[48][3]  ( .D(n7555), .CK(clk), .Q(\buff[48][3] ) );
  DFFQX1 \buff_reg[48][2]  ( .D(n2716), .CK(clk), .Q(\buff[48][2] ) );
  DFFQX1 \buff_reg[48][1]  ( .D(n2715), .CK(clk), .Q(\buff[48][1] ) );
  DFFQX1 \buff_reg[48][0]  ( .D(n7549), .CK(clk), .Q(\buff[48][0] ) );
  DFFQX1 \buff_reg[2][7]  ( .D(n7548), .CK(clk), .Q(\buff[2][7] ) );
  DFFQX1 \buff_reg[2][6]  ( .D(n7546), .CK(clk), .Q(\buff[2][6] ) );
  DFFQX1 \buff_reg[2][5]  ( .D(n8301), .CK(clk), .Q(\buff[2][5] ) );
  DFFQX1 \buff_reg[2][4]  ( .D(n8299), .CK(clk), .Q(\buff[2][4] ) );
  DFFQX1 \buff_reg[2][3]  ( .D(n8297), .CK(clk), .Q(\buff[2][3] ) );
  DFFQX1 \buff_reg[2][2]  ( .D(n8295), .CK(clk), .Q(\buff[2][2] ) );
  DFFQX1 \buff_reg[2][1]  ( .D(n8293), .CK(clk), .Q(\buff[2][1] ) );
  DFFQX1 \buff_reg[2][0]  ( .D(n8291), .CK(clk), .Q(\buff[2][0] ) );
  DFFQX1 \buff_reg[10][7]  ( .D(n3025), .CK(clk), .Q(\buff[10][7] ) );
  DFFQX1 \buff_reg[10][6]  ( .D(n3024), .CK(clk), .Q(\buff[10][6] ) );
  DFFQX1 \buff_reg[10][5]  ( .D(n3023), .CK(clk), .Q(\buff[10][5] ) );
  DFFQX1 \buff_reg[10][4]  ( .D(n3022), .CK(clk), .Q(\buff[10][4] ) );
  DFFQX1 \buff_reg[10][3]  ( .D(n3021), .CK(clk), .Q(\buff[10][3] ) );
  DFFQX1 \buff_reg[10][2]  ( .D(n3020), .CK(clk), .Q(\buff[10][2] ) );
  DFFQX1 \buff_reg[10][1]  ( .D(n3019), .CK(clk), .Q(\buff[10][1] ) );
  DFFQX1 \buff_reg[10][0]  ( .D(n8159), .CK(clk), .Q(\buff[10][0] ) );
  DFFQX1 \buff_reg[18][7]  ( .D(n2961), .CK(clk), .Q(\buff[18][7] ) );
  DFFQX1 \buff_reg[18][6]  ( .D(n2960), .CK(clk), .Q(\buff[18][6] ) );
  DFFQX1 \buff_reg[18][5]  ( .D(n2959), .CK(clk), .Q(\buff[18][5] ) );
  DFFQX1 \buff_reg[18][4]  ( .D(n2958), .CK(clk), .Q(\buff[18][4] ) );
  DFFQX1 \buff_reg[18][3]  ( .D(n2957), .CK(clk), .Q(\buff[18][3] ) );
  DFFQX1 \buff_reg[18][2]  ( .D(n2956), .CK(clk), .Q(\buff[18][2] ) );
  DFFQX1 \buff_reg[18][1]  ( .D(n2955), .CK(clk), .Q(\buff[18][1] ) );
  DFFQX1 \buff_reg[18][0]  ( .D(n8030), .CK(clk), .Q(\buff[18][0] ) );
  DFFQX1 \buff_reg[34][7]  ( .D(n8028), .CK(clk), .Q(\buff[34][7] ) );
  DFFQX1 \buff_reg[34][6]  ( .D(n8026), .CK(clk), .Q(\buff[34][6] ) );
  DFFQX1 \buff_reg[34][5]  ( .D(n2831), .CK(clk), .Q(\buff[34][5] ) );
  DFFQX1 \buff_reg[34][4]  ( .D(n2830), .CK(clk), .Q(\buff[34][4] ) );
  DFFQX1 \buff_reg[34][3]  ( .D(n2829), .CK(clk), .Q(\buff[34][3] ) );
  DFFQX1 \buff_reg[34][2]  ( .D(n2828), .CK(clk), .Q(\buff[34][2] ) );
  DFFQX1 \buff_reg[34][1]  ( .D(n7775), .CK(clk), .Q(\buff[34][1] ) );
  DFFQX1 \buff_reg[34][0]  ( .D(n7773), .CK(clk), .Q(\buff[34][0] ) );
  DFFQX1 \buff_reg[42][7]  ( .D(n2769), .CK(clk), .Q(\buff[42][7] ) );
  DFFQX1 \buff_reg[42][6]  ( .D(n2768), .CK(clk), .Q(\buff[42][6] ) );
  DFFQX1 \buff_reg[42][5]  ( .D(n2767), .CK(clk), .Q(\buff[42][5] ) );
  DFFQX1 \buff_reg[42][4]  ( .D(n2766), .CK(clk), .Q(\buff[42][4] ) );
  DFFQX1 \buff_reg[42][3]  ( .D(n2765), .CK(clk), .Q(\buff[42][3] ) );
  DFFQX1 \buff_reg[42][2]  ( .D(n2764), .CK(clk), .Q(\buff[42][2] ) );
  DFFQX1 \buff_reg[42][1]  ( .D(n2763), .CK(clk), .Q(\buff[42][1] ) );
  DFFQX1 \buff_reg[42][0]  ( .D(n7645), .CK(clk), .Q(\buff[42][0] ) );
  DFFQX1 \buff_reg[50][7]  ( .D(n7643), .CK(clk), .Q(\buff[50][7] ) );
  DFFQX1 \buff_reg[50][6]  ( .D(n7641), .CK(clk), .Q(\buff[50][6] ) );
  DFFQX1 \buff_reg[50][5]  ( .D(n7526), .CK(clk), .Q(\buff[50][5] ) );
  DFFQX1 \buff_reg[50][4]  ( .D(n7524), .CK(clk), .Q(\buff[50][4] ) );
  DFFQX1 \buff_reg[50][3]  ( .D(n2701), .CK(clk), .Q(\buff[50][3] ) );
  DFFQX1 \buff_reg[50][2]  ( .D(n2700), .CK(clk), .Q(\buff[50][2] ) );
  DFFQX1 \buff_reg[50][1]  ( .D(n2699), .CK(clk), .Q(\buff[50][1] ) );
  DFFQX1 \buff_reg[50][0]  ( .D(n7515), .CK(clk), .Q(\buff[50][0] ) );
  DFFQX1 \buff_reg[5][7]  ( .D(n3065), .CK(clk), .Q(\buff[5][7] ) );
  DFFQX1 \buff_reg[5][6]  ( .D(n3064), .CK(clk), .Q(\buff[5][6] ) );
  DFFQX1 \buff_reg[5][5]  ( .D(n8251), .CK(clk), .Q(\buff[5][5] ) );
  DFFQX1 \buff_reg[5][4]  ( .D(n3062), .CK(clk), .Q(\buff[5][4] ) );
  DFFQX1 \buff_reg[5][3]  ( .D(n8246), .CK(clk), .Q(\buff[5][3] ) );
  DFFQX1 \buff_reg[5][2]  ( .D(n8244), .CK(clk), .Q(\buff[5][2] ) );
  DFFQX1 \buff_reg[5][1]  ( .D(n8242), .CK(clk), .Q(\buff[5][1] ) );
  DFFQX1 \buff_reg[5][0]  ( .D(n8240), .CK(clk), .Q(\buff[5][0] ) );
  DFFQX1 \buff_reg[13][7]  ( .D(n8238), .CK(clk), .Q(\buff[13][7] ) );
  DFFQX1 \buff_reg[13][6]  ( .D(n8236), .CK(clk), .Q(\buff[13][6] ) );
  DFFQX1 \buff_reg[13][5]  ( .D(n2999), .CK(clk), .Q(\buff[13][5] ) );
  DFFQX1 \buff_reg[13][4]  ( .D(n2998), .CK(clk), .Q(\buff[13][4] ) );
  DFFQX1 \buff_reg[13][3]  ( .D(n2997), .CK(clk), .Q(\buff[13][3] ) );
  DFFQX1 \buff_reg[13][2]  ( .D(n2996), .CK(clk), .Q(\buff[13][2] ) );
  DFFQX1 \buff_reg[13][1]  ( .D(n2995), .CK(clk), .Q(\buff[13][1] ) );
  DFFQX1 \buff_reg[13][0]  ( .D(n8111), .CK(clk), .Q(\buff[13][0] ) );
  DFFQX1 \buff_reg[21][7]  ( .D(n8109), .CK(clk), .Q(\buff[21][7] ) );
  DFFQX1 \buff_reg[21][6]  ( .D(n2936), .CK(clk), .Q(\buff[21][6] ) );
  DFFQX1 \buff_reg[21][5]  ( .D(n7992), .CK(clk), .Q(\buff[21][5] ) );
  DFFQX1 \buff_reg[21][4]  ( .D(n7990), .CK(clk), .Q(\buff[21][4] ) );
  DFFQX1 \buff_reg[21][3]  ( .D(n7988), .CK(clk), .Q(\buff[21][3] ) );
  DFFQX1 \buff_reg[21][2]  ( .D(n7986), .CK(clk), .Q(\buff[21][2] ) );
  DFFQX1 \buff_reg[21][1]  ( .D(n7984), .CK(clk), .Q(\buff[21][1] ) );
  DFFQX1 \buff_reg[21][0]  ( .D(n7982), .CK(clk), .Q(\buff[21][0] ) );
  DFFQX1 \buff_reg[29][7]  ( .D(n2873), .CK(clk), .Q(\buff[29][7] ) );
  DFFQX1 \buff_reg[29][6]  ( .D(n2872), .CK(clk), .Q(\buff[29][6] ) );
  DFFQX1 \buff_reg[29][5]  ( .D(n7864), .CK(clk), .Q(\buff[29][5] ) );
  DFFQX1 \buff_reg[29][4]  ( .D(n7862), .CK(clk), .Q(\buff[29][4] ) );
  DFFQX1 \buff_reg[29][3]  ( .D(n7860), .CK(clk), .Q(\buff[29][3] ) );
  DFFQX1 \buff_reg[29][2]  ( .D(n7858), .CK(clk), .Q(\buff[29][2] ) );
  DFFQX1 \buff_reg[29][1]  ( .D(n7856), .CK(clk), .Q(\buff[29][1] ) );
  DFFQX1 \buff_reg[29][0]  ( .D(n7854), .CK(clk), .Q(\buff[29][0] ) );
  DFFQX1 \buff_reg[37][7]  ( .D(n7852), .CK(clk), .Q(\buff[37][7] ) );
  DFFQX1 \buff_reg[37][6]  ( .D(n7850), .CK(clk), .Q(\buff[37][6] ) );
  DFFQX1 \buff_reg[37][5]  ( .D(n7735), .CK(clk), .Q(\buff[37][5] ) );
  DFFQX1 \buff_reg[37][4]  ( .D(n7733), .CK(clk), .Q(\buff[37][4] ) );
  DFFQX1 \buff_reg[37][3]  ( .D(n7731), .CK(clk), .Q(\buff[37][3] ) );
  DFFQX1 \buff_reg[37][2]  ( .D(n7729), .CK(clk), .Q(\buff[37][2] ) );
  DFFQX1 \buff_reg[37][1]  ( .D(n7727), .CK(clk), .Q(\buff[37][1] ) );
  DFFQX1 \buff_reg[37][0]  ( .D(n7725), .CK(clk), .Q(\buff[37][0] ) );
  DFFQX1 \buff_reg[45][7]  ( .D(n2745), .CK(clk), .Q(\buff[45][7] ) );
  DFFQX1 \buff_reg[45][6]  ( .D(n2744), .CK(clk), .Q(\buff[45][6] ) );
  DFFQX1 \buff_reg[45][5]  ( .D(n7607), .CK(clk), .Q(\buff[45][5] ) );
  DFFQX1 \buff_reg[45][4]  ( .D(n7605), .CK(clk), .Q(\buff[45][4] ) );
  DFFQX1 \buff_reg[45][3]  ( .D(n7603), .CK(clk), .Q(\buff[45][3] ) );
  DFFQX1 \buff_reg[45][2]  ( .D(n7601), .CK(clk), .Q(\buff[45][2] ) );
  DFFQX1 \buff_reg[45][1]  ( .D(n7599), .CK(clk), .Q(\buff[45][1] ) );
  DFFQX1 \buff_reg[45][0]  ( .D(n7597), .CK(clk), .Q(\buff[45][0] ) );
  DFFQX1 \buff_reg[53][7]  ( .D(n7595), .CK(clk), .Q(\buff[53][7] ) );
  DFFQX1 \buff_reg[53][6]  ( .D(n7593), .CK(clk), .Q(\buff[53][6] ) );
  DFFQX1 \buff_reg[53][5]  ( .D(n7481), .CK(clk), .Q(\buff[53][5] ) );
  DFFQX1 \buff_reg[53][4]  ( .D(n7479), .CK(clk), .Q(\buff[53][4] ) );
  DFFQX1 \buff_reg[53][3]  ( .D(n7477), .CK(clk), .Q(\buff[53][3] ) );
  DFFQX1 \buff_reg[53][2]  ( .D(n2676), .CK(clk), .Q(\buff[53][2] ) );
  DFFQX1 \buff_reg[53][1]  ( .D(n7472), .CK(clk), .Q(\buff[53][1] ) );
  DFFQX1 \buff_reg[53][0]  ( .D(n7470), .CK(clk), .Q(\buff[53][0] ) );
  DFFQX1 \buff_reg[1][7]  ( .D(n3097), .CK(clk), .Q(\buff[1][7] ) );
  DFFQX1 \buff_reg[1][6]  ( .D(n3096), .CK(clk), .Q(\buff[1][6] ) );
  DFFQX1 \buff_reg[1][5]  ( .D(n8317), .CK(clk), .Q(\buff[1][5] ) );
  DFFQX1 \buff_reg[1][4]  ( .D(n8315), .CK(clk), .Q(\buff[1][4] ) );
  DFFQX1 \buff_reg[1][3]  ( .D(n3093), .CK(clk), .Q(\buff[1][3] ) );
  DFFQX1 \buff_reg[1][2]  ( .D(n8310), .CK(clk), .Q(\buff[1][2] ) );
  DFFQX1 \buff_reg[1][1]  ( .D(n8308), .CK(clk), .Q(\buff[1][1] ) );
  DFFQX1 \buff_reg[1][0]  ( .D(n8306), .CK(clk), .Q(\buff[1][0] ) );
  DFFQX1 \buff_reg[9][7]  ( .D(n3033), .CK(clk), .Q(\buff[9][7] ) );
  DFFQX1 \buff_reg[9][6]  ( .D(n3032), .CK(clk), .Q(\buff[9][6] ) );
  DFFQX1 \buff_reg[9][5]  ( .D(n8185), .CK(clk), .Q(\buff[9][5] ) );
  DFFQX1 \buff_reg[9][4]  ( .D(n8183), .CK(clk), .Q(\buff[9][4] ) );
  DFFQX1 \buff_reg[9][3]  ( .D(n8181), .CK(clk), .Q(\buff[9][3] ) );
  DFFQX1 \buff_reg[9][2]  ( .D(n8179), .CK(clk), .Q(\buff[9][2] ) );
  DFFQX1 \buff_reg[9][1]  ( .D(n8177), .CK(clk), .Q(\buff[9][1] ) );
  DFFQX1 \buff_reg[9][0]  ( .D(n8175), .CK(clk), .Q(\buff[9][0] ) );
  DFFQX1 \buff_reg[17][7]  ( .D(n2969), .CK(clk), .Q(\buff[17][7] ) );
  DFFQX1 \buff_reg[17][6]  ( .D(n2968), .CK(clk), .Q(\buff[17][6] ) );
  DFFQX1 \buff_reg[17][5]  ( .D(n8056), .CK(clk), .Q(\buff[17][5] ) );
  DFFQX1 \buff_reg[17][4]  ( .D(n8054), .CK(clk), .Q(\buff[17][4] ) );
  DFFQX1 \buff_reg[17][3]  ( .D(n8052), .CK(clk), .Q(\buff[17][3] ) );
  DFFQX1 \buff_reg[17][2]  ( .D(n8050), .CK(clk), .Q(\buff[17][2] ) );
  DFFQX1 \buff_reg[17][1]  ( .D(n8048), .CK(clk), .Q(\buff[17][1] ) );
  DFFQX1 \buff_reg[17][0]  ( .D(n8046), .CK(clk), .Q(\buff[17][0] ) );
  DFFQX1 \buff_reg[25][7]  ( .D(n2905), .CK(clk), .Q(\buff[25][7] ) );
  DFFQX1 \buff_reg[25][6]  ( .D(n2904), .CK(clk), .Q(\buff[25][6] ) );
  DFFQX1 \buff_reg[25][5]  ( .D(n7928), .CK(clk), .Q(\buff[25][5] ) );
  DFFQX1 \buff_reg[25][4]  ( .D(n7926), .CK(clk), .Q(\buff[25][4] ) );
  DFFQX1 \buff_reg[25][3]  ( .D(n7924), .CK(clk), .Q(\buff[25][3] ) );
  DFFQX1 \buff_reg[25][2]  ( .D(n7922), .CK(clk), .Q(\buff[25][2] ) );
  DFFQX1 \buff_reg[25][1]  ( .D(n7920), .CK(clk), .Q(\buff[25][1] ) );
  DFFQX1 \buff_reg[25][0]  ( .D(n7918), .CK(clk), .Q(\buff[25][0] ) );
  DFFQX1 \buff_reg[33][7]  ( .D(n7916), .CK(clk), .Q(\buff[33][7] ) );
  DFFQX1 \buff_reg[33][6]  ( .D(n7914), .CK(clk), .Q(\buff[33][6] ) );
  DFFQX1 \buff_reg[33][5]  ( .D(n7799), .CK(clk), .Q(\buff[33][5] ) );
  DFFQX1 \buff_reg[33][4]  ( .D(n7797), .CK(clk), .Q(\buff[33][4] ) );
  DFFQX1 \buff_reg[33][3]  ( .D(n7795), .CK(clk), .Q(\buff[33][3] ) );
  DFFQX1 \buff_reg[33][2]  ( .D(n7793), .CK(clk), .Q(\buff[33][2] ) );
  DFFQX1 \buff_reg[33][1]  ( .D(n7791), .CK(clk), .Q(\buff[33][1] ) );
  DFFQX1 \buff_reg[33][0]  ( .D(n7789), .CK(clk), .Q(\buff[33][0] ) );
  DFFQX1 \buff_reg[41][7]  ( .D(n2777), .CK(clk), .Q(\buff[41][7] ) );
  DFFQX1 \buff_reg[41][6]  ( .D(n2776), .CK(clk), .Q(\buff[41][6] ) );
  DFFQX1 \buff_reg[41][5]  ( .D(n7671), .CK(clk), .Q(\buff[41][5] ) );
  DFFQX1 \buff_reg[41][4]  ( .D(n7669), .CK(clk), .Q(\buff[41][4] ) );
  DFFQX1 \buff_reg[41][3]  ( .D(n7667), .CK(clk), .Q(\buff[41][3] ) );
  DFFQX1 \buff_reg[41][2]  ( .D(n7665), .CK(clk), .Q(\buff[41][2] ) );
  DFFQX1 \buff_reg[41][1]  ( .D(n7663), .CK(clk), .Q(\buff[41][1] ) );
  DFFQX1 \buff_reg[41][0]  ( .D(n7661), .CK(clk), .Q(\buff[41][0] ) );
  DFFQX1 \buff_reg[49][7]  ( .D(n7659), .CK(clk), .Q(\buff[49][7] ) );
  DFFQX1 \buff_reg[49][6]  ( .D(n7657), .CK(clk), .Q(\buff[49][6] ) );
  DFFQX1 \buff_reg[49][5]  ( .D(n7543), .CK(clk), .Q(\buff[49][5] ) );
  DFFQX1 \buff_reg[49][4]  ( .D(n7541), .CK(clk), .Q(\buff[49][4] ) );
  DFFQX1 \buff_reg[49][3]  ( .D(n2709), .CK(clk), .Q(\buff[49][3] ) );
  DFFQX1 \buff_reg[49][2]  ( .D(n7536), .CK(clk), .Q(\buff[49][2] ) );
  DFFQX1 \buff_reg[49][1]  ( .D(n7534), .CK(clk), .Q(\buff[49][1] ) );
  DFFQX1 \buff_reg[49][0]  ( .D(n7532), .CK(clk), .Q(\buff[49][0] ) );
  DFFQX1 \buff_reg[55][7]  ( .D(n2665), .CK(clk), .Q(\buff[55][7] ) );
  DFFQX1 \buff_reg[55][6]  ( .D(n2664), .CK(clk), .Q(\buff[55][6] ) );
  DFFQX1 \buff_reg[55][5]  ( .D(n2663), .CK(clk), .Q(\buff[55][5] ) );
  DFFQX1 \buff_reg[55][4]  ( .D(n7447), .CK(clk), .Q(\buff[55][4] ) );
  DFFQX1 \buff_reg[55][3]  ( .D(n7444), .CK(clk), .Q(\buff[55][3] ) );
  DFFQX1 \buff_reg[55][2]  ( .D(n7442), .CK(clk), .Q(\buff[55][2] ) );
  DFFQX1 \buff_reg[55][1]  ( .D(n7440), .CK(clk), .Q(\buff[55][1] ) );
  DFFQX1 \buff_reg[55][0]  ( .D(n7438), .CK(clk), .Q(\buff[55][0] ) );
  DFFQX1 \buff_reg[23][7]  ( .D(n7437), .CK(clk), .Q(\buff[23][7] ) );
  DFFQX1 \buff_reg[23][6]  ( .D(n8354), .CK(clk), .Q(\buff[23][6] ) );
  DFFQX1 \buff_reg[23][5]  ( .D(n7961), .CK(clk), .Q(\buff[23][5] ) );
  DFFQX1 \buff_reg[23][4]  ( .D(n7958), .CK(clk), .Q(\buff[23][4] ) );
  DFFQX1 \buff_reg[23][3]  ( .D(n7956), .CK(clk), .Q(\buff[23][3] ) );
  DFFQX1 \buff_reg[23][2]  ( .D(n7954), .CK(clk), .Q(\buff[23][2] ) );
  DFFQX1 \buff_reg[23][1]  ( .D(n7952), .CK(clk), .Q(\buff[23][1] ) );
  DFFQX1 \buff_reg[23][0]  ( .D(n7950), .CK(clk), .Q(\buff[23][0] ) );
  DFFQX1 \buff_reg[27][7]  ( .D(n7949), .CK(clk), .Q(\buff[27][7] ) );
  DFFQX1 \buff_reg[27][6]  ( .D(n2888), .CK(clk), .Q(\buff[27][6] ) );
  DFFQX1 \buff_reg[27][5]  ( .D(n7897), .CK(clk), .Q(\buff[27][5] ) );
  DFFQX1 \buff_reg[27][4]  ( .D(n7895), .CK(clk), .Q(\buff[27][4] ) );
  DFFQX1 \buff_reg[27][3]  ( .D(n7893), .CK(clk), .Q(\buff[27][3] ) );
  DFFQX1 \buff_reg[27][2]  ( .D(n7891), .CK(clk), .Q(\buff[27][2] ) );
  DFFQX1 \buff_reg[27][1]  ( .D(n7889), .CK(clk), .Q(\buff[27][1] ) );
  DFFQX1 \buff_reg[27][0]  ( .D(n7887), .CK(clk), .Q(\buff[27][0] ) );
  DFFRX1 \cnt_reg[6]  ( .D(n7499), .CK(clk), .RN(n9669), .Q(\cnt[6] ), .QN(
        n2581) );
  DFFQX1 \buff_reg[7][7]  ( .D(n8353), .CK(clk), .Q(\buff[7][7] ) );
  DFFQX1 \buff_reg[7][6]  ( .D(n8341), .CK(clk), .Q(\buff[7][6] ) );
  DFFQX1 \buff_reg[7][5]  ( .D(n7885), .CK(clk), .Q(\buff[7][5] ) );
  DFFQX1 \buff_reg[7][4]  ( .D(n7882), .CK(clk), .Q(\buff[7][4] ) );
  DFFQX1 \buff_reg[7][3]  ( .D(n8218), .CK(clk), .Q(\buff[7][3] ) );
  DFFQX1 \buff_reg[7][2]  ( .D(n8216), .CK(clk), .Q(\buff[7][2] ) );
  DFFQX1 \buff_reg[7][1]  ( .D(n8214), .CK(clk), .Q(\buff[7][1] ) );
  DFFQX1 \buff_reg[7][0]  ( .D(n8212), .CK(clk), .Q(\buff[7][0] ) );
  DFFQX1 \buff_reg[15][7]  ( .D(n8211), .CK(clk), .Q(\buff[15][7] ) );
  DFFQX1 \buff_reg[15][6]  ( .D(n8209), .CK(clk), .Q(\buff[15][6] ) );
  DFFQX1 \buff_reg[15][5]  ( .D(n8207), .CK(clk), .Q(\buff[15][5] ) );
  DFFQX1 \buff_reg[15][4]  ( .D(n8205), .CK(clk), .Q(\buff[15][4] ) );
  DFFQX1 \buff_reg[15][3]  ( .D(n8088), .CK(clk), .Q(\buff[15][3] ) );
  DFFQX1 \buff_reg[15][2]  ( .D(n8086), .CK(clk), .Q(\buff[15][2] ) );
  DFFQX1 \buff_reg[15][1]  ( .D(n8084), .CK(clk), .Q(\buff[15][1] ) );
  DFFQX1 \buff_reg[15][0]  ( .D(n8082), .CK(clk), .Q(\buff[15][0] ) );
  DFFQX1 \buff_reg[31][7]  ( .D(n8081), .CK(clk), .Q(\buff[31][7] ) );
  DFFQX1 \buff_reg[31][6]  ( .D(n8078), .CK(clk), .Q(\buff[31][6] ) );
  DFFQX1 \buff_reg[31][5]  ( .D(n8077), .CK(clk), .Q(\buff[31][5] ) );
  DFFQX1 \buff_reg[31][4]  ( .D(n8075), .CK(clk), .Q(\buff[31][4] ) );
  DFFQX1 \buff_reg[31][3]  ( .D(n7833), .CK(clk), .Q(\buff[31][3] ) );
  DFFQX1 \buff_reg[31][2]  ( .D(n7831), .CK(clk), .Q(\buff[31][2] ) );
  DFFQX1 \buff_reg[31][1]  ( .D(n7829), .CK(clk), .Q(\buff[31][1] ) );
  DFFQX1 \buff_reg[31][0]  ( .D(n7826), .CK(clk), .Q(\buff[31][0] ) );
  DFFQX1 \buff_reg[39][7]  ( .D(n7825), .CK(clk), .Q(\buff[39][7] ) );
  DFFQX1 \buff_reg[39][6]  ( .D(n7822), .CK(clk), .Q(\buff[39][6] ) );
  DFFQX1 \buff_reg[39][5]  ( .D(n7821), .CK(clk), .Q(\buff[39][5] ) );
  DFFQX1 \buff_reg[39][4]  ( .D(n7819), .CK(clk), .Q(\buff[39][4] ) );
  DFFQX1 \buff_reg[39][3]  ( .D(n7704), .CK(clk), .Q(\buff[39][3] ) );
  DFFQX1 \buff_reg[39][2]  ( .D(n7702), .CK(clk), .Q(\buff[39][2] ) );
  DFFQX1 \buff_reg[39][1]  ( .D(n7700), .CK(clk), .Q(\buff[39][1] ) );
  DFFQX1 \buff_reg[39][0]  ( .D(n7697), .CK(clk), .Q(\buff[39][0] ) );
  DFFQX1 \buff_reg[47][7]  ( .D(n7696), .CK(clk), .Q(\buff[47][7] ) );
  DFFQX1 \buff_reg[47][6]  ( .D(n7693), .CK(clk), .Q(\buff[47][6] ) );
  DFFQX1 \buff_reg[47][5]  ( .D(n7692), .CK(clk), .Q(\buff[47][5] ) );
  DFFQX1 \buff_reg[47][4]  ( .D(n7690), .CK(clk), .Q(\buff[47][4] ) );
  DFFQX1 \buff_reg[47][3]  ( .D(n7576), .CK(clk), .Q(\buff[47][3] ) );
  DFFQX1 \buff_reg[47][2]  ( .D(n7574), .CK(clk), .Q(\buff[47][2] ) );
  DFFQX1 \buff_reg[47][1]  ( .D(n7572), .CK(clk), .Q(\buff[47][1] ) );
  DFFQX1 \buff_reg[47][0]  ( .D(n7569), .CK(clk), .Q(\buff[47][0] ) );
  DFFQX1 \buff_reg[3][7]  ( .D(n7567), .CK(clk), .Q(\buff[3][7] ) );
  DFFQX1 \buff_reg[3][6]  ( .D(n7565), .CK(clk), .Q(\buff[3][6] ) );
  DFFQX1 \buff_reg[3][5]  ( .D(n7563), .CK(clk), .Q(\buff[3][5] ) );
  DFFQX1 \buff_reg[3][4]  ( .D(n7561), .CK(clk), .Q(\buff[3][4] ) );
  DFFQX1 \buff_reg[3][3]  ( .D(n8284), .CK(clk), .Q(\buff[3][3] ) );
  DFFQX1 \buff_reg[3][2]  ( .D(n8282), .CK(clk), .Q(\buff[3][2] ) );
  DFFQX1 \buff_reg[3][1]  ( .D(n8280), .CK(clk), .Q(\buff[3][1] ) );
  DFFQX1 \buff_reg[3][0]  ( .D(n8278), .CK(clk), .Q(\buff[3][0] ) );
  DFFQX1 \buff_reg[11][7]  ( .D(n8276), .CK(clk), .Q(\buff[11][7] ) );
  DFFQX1 \buff_reg[11][6]  ( .D(n8274), .CK(clk), .Q(\buff[11][6] ) );
  DFFQX1 \buff_reg[11][5]  ( .D(n8272), .CK(clk), .Q(\buff[11][5] ) );
  DFFQX1 \buff_reg[11][4]  ( .D(n8270), .CK(clk), .Q(\buff[11][4] ) );
  DFFQX1 \buff_reg[11][3]  ( .D(n8153), .CK(clk), .Q(\buff[11][3] ) );
  DFFQX1 \buff_reg[11][2]  ( .D(n8151), .CK(clk), .Q(\buff[11][2] ) );
  DFFQX1 \buff_reg[11][1]  ( .D(n8149), .CK(clk), .Q(\buff[11][1] ) );
  DFFQX1 \buff_reg[11][0]  ( .D(n8147), .CK(clk), .Q(\buff[11][0] ) );
  DFFQX1 \buff_reg[19][7]  ( .D(n8145), .CK(clk), .Q(\buff[19][7] ) );
  DFFQX1 \buff_reg[19][6]  ( .D(n8143), .CK(clk), .Q(\buff[19][6] ) );
  DFFQX1 \buff_reg[19][5]  ( .D(n8141), .CK(clk), .Q(\buff[19][5] ) );
  DFFQX1 \buff_reg[19][4]  ( .D(n8139), .CK(clk), .Q(\buff[19][4] ) );
  DFFQX1 \buff_reg[19][3]  ( .D(n8024), .CK(clk), .Q(\buff[19][3] ) );
  DFFQX1 \buff_reg[19][2]  ( .D(n8022), .CK(clk), .Q(\buff[19][2] ) );
  DFFQX1 \buff_reg[19][1]  ( .D(n8020), .CK(clk), .Q(\buff[19][1] ) );
  DFFQX1 \buff_reg[19][0]  ( .D(n8018), .CK(clk), .Q(\buff[19][0] ) );
  DFFQX1 \buff_reg[35][7]  ( .D(n8016), .CK(clk), .Q(\buff[35][7] ) );
  DFFQX1 \buff_reg[35][6]  ( .D(n8014), .CK(clk), .Q(\buff[35][6] ) );
  DFFQX1 \buff_reg[35][5]  ( .D(n8012), .CK(clk), .Q(\buff[35][5] ) );
  DFFQX1 \buff_reg[35][4]  ( .D(n8010), .CK(clk), .Q(\buff[35][4] ) );
  DFFQX1 \buff_reg[35][3]  ( .D(n7767), .CK(clk), .Q(\buff[35][3] ) );
  DFFQX1 \buff_reg[35][2]  ( .D(n7765), .CK(clk), .Q(\buff[35][2] ) );
  DFFQX1 \buff_reg[35][1]  ( .D(n7763), .CK(clk), .Q(\buff[35][1] ) );
  DFFQX1 \buff_reg[35][0]  ( .D(n7761), .CK(clk), .Q(\buff[35][0] ) );
  DFFQX1 \buff_reg[43][7]  ( .D(n7759), .CK(clk), .Q(\buff[43][7] ) );
  DFFQX1 \buff_reg[43][6]  ( .D(n7757), .CK(clk), .Q(\buff[43][6] ) );
  DFFQX1 \buff_reg[43][5]  ( .D(n7755), .CK(clk), .Q(\buff[43][5] ) );
  DFFQX1 \buff_reg[43][4]  ( .D(n7753), .CK(clk), .Q(\buff[43][4] ) );
  DFFQX1 \buff_reg[43][3]  ( .D(n7639), .CK(clk), .Q(\buff[43][3] ) );
  DFFQX1 \buff_reg[43][2]  ( .D(n7637), .CK(clk), .Q(\buff[43][2] ) );
  DFFQX1 \buff_reg[43][1]  ( .D(n7635), .CK(clk), .Q(\buff[43][1] ) );
  DFFQX1 \buff_reg[43][0]  ( .D(n7633), .CK(clk), .Q(\buff[43][0] ) );
  DFFQX1 \buff_reg[51][7]  ( .D(n7631), .CK(clk), .Q(\buff[51][7] ) );
  DFFQX1 \buff_reg[51][6]  ( .D(n7629), .CK(clk), .Q(\buff[51][6] ) );
  DFFQX1 \buff_reg[51][5]  ( .D(n7627), .CK(clk), .Q(\buff[51][5] ) );
  DFFQX1 \buff_reg[51][4]  ( .D(n7625), .CK(clk), .Q(\buff[51][4] ) );
  DFFQX1 \buff_reg[51][3]  ( .D(n7509), .CK(clk), .Q(\buff[51][3] ) );
  DFFQX1 \buff_reg[51][2]  ( .D(n7507), .CK(clk), .Q(\buff[51][2] ) );
  DFFQX1 \buff_reg[51][1]  ( .D(n7505), .CK(clk), .Q(\buff[51][1] ) );
  DFFQX1 \buff_reg[51][0]  ( .D(n7503), .CK(clk), .Q(\buff[51][0] ) );
  DFFSX4 \x_reg[2]  ( .D(n8364), .CK(clk), .SN(n9669), .Q(n8431), .QN(n2575)
         );
  DFFRX1 \x_reg[1]  ( .D(n8359), .CK(clk), .RN(n9459), .Q(n8416), .QN(n2576)
         );
  DFFRX1 IROM_EN_reg ( .D(n8351), .CK(clk), .RN(n9459), .Q(n9830), .QN(n2572)
         );
  DFFSX1 busy_reg ( .D(n8339), .CK(clk), .SN(n9669), .Q(n9846), .QN(n2588) );
  DFFRX1 \cnt_reg[2]  ( .D(n8343), .CK(clk), .RN(n9669), .Q(N1658), .QN(n2585)
         );
  DFFSRXL \cur_reg[1]  ( .D(n8345), .CK(clk), .SN(1'b1), .RN(n9669), .QN(n2571) );
  DFFSRXL \cur_reg[0]  ( .D(n8347), .CK(clk), .SN(1'b1), .RN(n9669), .Q(n9743), 
        .QN(n2574) );
  DFFSX1 \y_reg[2]  ( .D(n7501), .CK(clk), .SN(n9669), .Q(n9515), .QN(n9514)
         );
  EDFFX1 \cmd_reg_reg[2]  ( .D(cmd[2]), .E(n2593), .CK(clk), .Q(n9747), .QN(
        n2589) );
  EDFFX1 \cmd_reg_reg[1]  ( .D(cmd[1]), .E(n2593), .CK(clk), .Q(n9748), .QN(
        n2590) );
  EDFFX1 \cmd_reg_reg[0]  ( .D(cmd[0]), .E(n2593), .CK(clk), .Q(n9738), .QN(
        n2591) );
  DFFRX4 \cnt_reg[5]  ( .D(n8386), .CK(clk), .RN(n9669), .Q(N1661), .QN(n2582)
         );
  DFFRX2 \cnt_reg[3]  ( .D(n8374), .CK(clk), .RN(n9669), .Q(N1659), .QN(n2584)
         );
  DFFRX2 \cnt_reg[1]  ( .D(n8376), .CK(clk), .RN(n9669), .Q(N1657), .QN(n2586)
         );
  DFFRX2 \cnt_reg[0]  ( .D(n8379), .CK(clk), .RN(n9669), .Q(N1656), .QN(n2587)
         );
  DFFSRX2 \x_reg[0]  ( .D(n8371), .CK(clk), .SN(1'b1), .RN(n9669), .Q(n9517), 
        .QN(n9516) );
  DFFSRX2 \y_reg[0]  ( .D(n8369), .CK(clk), .SN(1'b1), .RN(n9669), .Q(n9511), 
        .QN(n9510) );
  DFFSRX2 \y_reg[1]  ( .D(n8366), .CK(clk), .SN(1'b1), .RN(n9669), .Q(n9513), 
        .QN(n9512) );
  DFFRX1 \cnt_reg[4]  ( .D(n8382), .CK(clk), .RN(n9669), .QN(n2583) );
  CLKBUFX2 U7143 ( .A(n2289), .Y(n9340) );
  NAND2X1 U7144 ( .A(n9662), .B(n2011), .Y(n1977) );
  BUFX2 U7145 ( .A(n1977), .Y(n7224) );
  CLKBUFX2 U7146 ( .A(n9517), .Y(n8373) );
  XNOR2XL U7147 ( .A(n2549), .B(n8373), .Y(n3110) );
  CLKBUFX8 U7148 ( .A(n280), .Y(n7225) );
  CLKBUFX8 U7149 ( .A(n259), .Y(n7226) );
  CLKINVX1 U7150 ( .A(n8740), .Y(n8903) );
  CLKINVX1 U7151 ( .A(n8747), .Y(n8904) );
  CLKINVX1 U7152 ( .A(\buff[11][2] ), .Y(n8865) );
  CLKINVX1 U7153 ( .A(n8754), .Y(n8905) );
  CLKINVX1 U7154 ( .A(n8761), .Y(n8906) );
  CLKINVX1 U7155 ( .A(\buff[11][5] ), .Y(n8868) );
  CLKINVX1 U7156 ( .A(n8775), .Y(n8908) );
  CLKINVX1 U7157 ( .A(n8782), .Y(n8909) );
  CLKINVX1 U7158 ( .A(n8789), .Y(n8910) );
  MXI3XL U7159 ( .A(n8491), .B(n8492), .C(n8493), .S0(n9513), .S1(n8928), .Y(
        n8490) );
  MXI3X1 U7160 ( .A(n8511), .B(n8512), .C(n8513), .S0(n9137), .S1(n8928), .Y(
        n8510) );
  MXI3X1 U7161 ( .A(n8571), .B(n8572), .C(n8573), .S0(n8924), .S1(n8928), .Y(
        n8570) );
  CLKINVX1 U7162 ( .A(\buff[11][0] ), .Y(n8863) );
  CLKINVX1 U7163 ( .A(\buff[11][3] ), .Y(n8866) );
  CLKINVX1 U7164 ( .A(\buff[11][4] ), .Y(n8867) );
  CLKINVX1 U7165 ( .A(\buff[11][6] ), .Y(n8869) );
  CLKINVX1 U7166 ( .A(\buff[7][7] ), .Y(n8878) );
  CLKBUFX3 U7167 ( .A(n160), .Y(n8106) );
  INVX3 U7168 ( .A(n9613), .Y(n9615) );
  INVX1 U7169 ( .A(n8794), .Y(N7388) );
  AOI2BB2X2 U7170 ( .B0(n9608), .B1(n9755), .A0N(n9615), .A1N(n9533), .Y(n626)
         );
  AOI2BB2X2 U7171 ( .B0(n9610), .B1(n9780), .A0N(n9615), .A1N(n9531), .Y(n950)
         );
  AOI2BB2X2 U7172 ( .B0(n9609), .B1(n9761), .A0N(n9615), .A1N(n9527), .Y(n1270) );
  NAND3X1 U7173 ( .A(n2584), .B(n8393), .C(n8385), .Y(n1654) );
  AOI2BB2X2 U7174 ( .B0(n9608), .B1(n9773), .A0N(n9614), .A1N(n7236), .Y(n2221) );
  AOI2BB2X2 U7175 ( .B0(n9609), .B1(n9758), .A0N(n9615), .A1N(n9387), .Y(n1428) );
  AOI2BB2X2 U7176 ( .B0(n9609), .B1(n9788), .A0N(n9614), .A1N(n9525), .Y(n1587) );
  CLKINVX1 U7177 ( .A(\buff[7][1] ), .Y(n8872) );
  CLKINVX1 U7178 ( .A(n8768), .Y(n8907) );
  OAI22XL U7179 ( .A0(n8312), .A1(n365), .B0(n367), .B1(n572), .Y(n571) );
  OAI22XL U7180 ( .A0(n9340), .A1(n160), .B0(n412), .B1(n2290), .Y(n2331) );
  OAI22XL U7181 ( .A0(n199), .A1(n365), .B0(n367), .B1(n532), .Y(n531) );
  AOI2BB2X2 U7182 ( .B0(n9608), .B1(n9769), .A0N(n9614), .A1N(n9361), .Y(n2422) );
  AOI2BB2X2 U7183 ( .B0(n9608), .B1(n9767), .A0N(n9614), .A1N(n9371), .Y(n1941) );
  NAND3X1 U7184 ( .A(n2587), .B(N1657), .C(n2132), .Y(n212) );
  MXI3X1 U7185 ( .A(n8531), .B(n8532), .C(n8533), .S0(n9137), .S1(n8928), .Y(
        n8530) );
  MXI3X1 U7186 ( .A(n8551), .B(n8552), .C(n8553), .S0(n8927), .S1(n8928), .Y(
        n8550) );
  MXI3X1 U7187 ( .A(n8591), .B(n8592), .C(n8593), .S0(n8924), .S1(n8928), .Y(
        n8590) );
  MXI3X1 U7188 ( .A(n8611), .B(n8612), .C(n8613), .S0(n8925), .S1(n8928), .Y(
        n8610) );
  MXI3X1 U7189 ( .A(n8631), .B(n8632), .C(n8633), .S0(n8925), .S1(n8928), .Y(
        n8630) );
  NAND2X1 U7190 ( .A(n9663), .B(n571), .Y(n537) );
  DLY4X1 U7191 ( .A(\buff[59][5] ), .Y(n7365) );
  DLY4X1 U7192 ( .A(\buff[59][7] ), .Y(n7299) );
  OA22X1 U7193 ( .A0(n159), .A1(n160), .B0(n161), .B1(n145), .Y(n148) );
  DLY4X1 U7194 ( .A(\buff[63][5] ), .Y(n7269) );
  DLY4X1 U7195 ( .A(\buff[63][6] ), .Y(n8363) );
  CLKBUFX3 U7196 ( .A(n119), .Y(n9438) );
  DLY4X1 U7197 ( .A(\buff[63][7] ), .Y(n8338) );
  DLY4X1 U7198 ( .A(n3114), .Y(n8384) );
  XNOR2X1 U7199 ( .A(n2538), .B(n8370), .Y(n3107) );
  CLKBUFX3 U7200 ( .A(next[1]), .Y(n8346) );
  OAI2BB2XL U7201 ( .B0(IRB_RW), .B1(n91), .A0N(n92), .A1N(n9663), .Y(next[1])
         );
  DLY4X1 U7202 ( .A(n3116), .Y(n8344) );
  DLY4X1 U7203 ( .A(n2573), .Y(n8351) );
  DLY4X1 U7204 ( .A(n3109), .Y(n8360) );
  OAI31XL U7205 ( .A0(n2549), .A1(n9813), .A2(n9737), .B0(n2555), .Y(n3111) );
  DLY3X1 U7206 ( .A(n2722), .Y(n7570) );
  DLY4X1 U7207 ( .A(n2723), .Y(n7572) );
  DLY4X1 U7208 ( .A(n2724), .Y(n7574) );
  DLY4X1 U7209 ( .A(n2725), .Y(n7576) );
  DLY4X1 U7210 ( .A(n2726), .Y(n7690) );
  DLY4X1 U7211 ( .A(n2727), .Y(n7692) );
  DLY3X1 U7212 ( .A(n2786), .Y(n7698) );
  DLY4X1 U7213 ( .A(n2787), .Y(n7700) );
  DLY4X1 U7214 ( .A(n2788), .Y(n7702) );
  DLY4X1 U7215 ( .A(n2789), .Y(n7704) );
  DLY4X1 U7216 ( .A(n2790), .Y(n7819) );
  DLY4X1 U7217 ( .A(n2791), .Y(n7821) );
  DLY3X1 U7218 ( .A(n2850), .Y(n7827) );
  DLY4X1 U7219 ( .A(n2851), .Y(n7829) );
  DLY4X1 U7220 ( .A(n2852), .Y(n7831) );
  DLY4X1 U7221 ( .A(n2853), .Y(n7833) );
  DLY4X1 U7222 ( .A(n2854), .Y(n8075) );
  DLY4X1 U7223 ( .A(n2855), .Y(n8077) );
  DLY4X1 U7224 ( .A(n2857), .Y(n8081) );
  DLY3X1 U7225 ( .A(n2978), .Y(n8083) );
  DLY3X1 U7226 ( .A(n2979), .Y(n8085) );
  DLY3X1 U7227 ( .A(n2980), .Y(n8087) );
  DLY3X1 U7228 ( .A(n2981), .Y(n8089) );
  DLY4X1 U7229 ( .A(n2982), .Y(n8205) );
  DLY4X1 U7230 ( .A(n2983), .Y(n8207) );
  DLY4X1 U7231 ( .A(n2984), .Y(n8209) );
  DLY4X1 U7232 ( .A(n2985), .Y(n8211) );
  DLY3X1 U7233 ( .A(n3042), .Y(n8213) );
  DLY3X1 U7234 ( .A(n3043), .Y(n8215) );
  DLY3X1 U7235 ( .A(n3044), .Y(n8217) );
  DLY3X1 U7236 ( .A(n3045), .Y(n8219) );
  DLY3X1 U7237 ( .A(n3046), .Y(n7883) );
  DLY4X1 U7238 ( .A(n3119), .Y(n7500) );
  DLY4X1 U7239 ( .A(n2882), .Y(n7887) );
  DLY4X1 U7240 ( .A(n2883), .Y(n7889) );
  DLY4X1 U7241 ( .A(n2884), .Y(n7891) );
  DLY4X1 U7242 ( .A(n2885), .Y(n7893) );
  DLY4X1 U7243 ( .A(n2886), .Y(n7895) );
  DLY4X1 U7244 ( .A(n2887), .Y(n7897) );
  DLY4X1 U7245 ( .A(n2889), .Y(n7949) );
  DLY4X1 U7246 ( .A(n2914), .Y(n7951) );
  DLY4X1 U7247 ( .A(n2915), .Y(n7953) );
  DLY4X1 U7248 ( .A(n2916), .Y(n7955) );
  DLY4X1 U7249 ( .A(n2917), .Y(n7957) );
  DLY4X1 U7250 ( .A(n2918), .Y(n7959) );
  DLY4X1 U7251 ( .A(n2658), .Y(n7439) );
  DLY4X1 U7252 ( .A(n2659), .Y(n7441) );
  DLY4X1 U7253 ( .A(n3082), .Y(n8291) );
  DLY4X1 U7254 ( .A(n3083), .Y(n8293) );
  DLY4X1 U7255 ( .A(n3084), .Y(n8295) );
  DLY4X1 U7256 ( .A(n3085), .Y(n8297) );
  DLY4X1 U7257 ( .A(n3086), .Y(n8299) );
  DLY4X1 U7258 ( .A(n3087), .Y(n8301) );
  DLY4X1 U7259 ( .A(n3089), .Y(n7548) );
  DLY4X1 U7260 ( .A(n2986), .Y(n8095) );
  DLY4X1 U7261 ( .A(n2987), .Y(n8097) );
  DLY4X1 U7262 ( .A(n2988), .Y(n8099) );
  DLY4X1 U7263 ( .A(n2989), .Y(n8101) );
  DLY4X1 U7264 ( .A(n2990), .Y(n8103) );
  DLY4X1 U7265 ( .A(n2630), .Y(n7362) );
  CLKMX2X2 U7266 ( .A(n8440), .B(n8672), .S0(n8919), .Y(n7227) );
  CLKMX2X2 U7267 ( .A(n8446), .B(n8698), .S0(n9125), .Y(n7228) );
  CLKMX2X2 U7268 ( .A(n8447), .B(n8711), .S0(n9126), .Y(n7229) );
  CLKMX2X2 U7269 ( .A(n8448), .B(n8724), .S0(n9126), .Y(n7230) );
  CLKMX2X2 U7270 ( .A(n8449), .B(n8737), .S0(n9129), .Y(n7231) );
  AOI22X1 U7271 ( .A0(n9617), .A1(N7395), .B0(n9607), .B1(n7231), .Y(n7232) );
  MX4X1 U7272 ( .A(n8913), .B(n8423), .C(n8757), .D(n8753), .S0(n9129), .S1(
        n8929), .Y(n7233) );
  CLKMX2X2 U7273 ( .A(n8441), .B(n8685), .S0(n8919), .Y(n7234) );
  MX4X1 U7274 ( .A(n8917), .B(n8427), .C(n8785), .D(n8781), .S0(n9129), .S1(
        n8929), .Y(n7235) );
  CLKBUFX2 U7275 ( .A(n9666), .Y(n9664) );
  NAND2X4 U7276 ( .A(n2211), .B(n667), .Y(n7236) );
  AOI22X1 U7277 ( .A0(n292), .A1(N7392), .B0(n9607), .B1(n7228), .Y(n7237) );
  AOI22X1 U7278 ( .A0(n9617), .A1(n7235), .B0(n9607), .B1(n7230), .Y(n7238) );
  AOI22X1 U7279 ( .A0(n9613), .A1(N7391), .B0(n9608), .B1(n7234), .Y(n7239) );
  AOI22X1 U7280 ( .A0(n292), .A1(n7233), .B0(n9607), .B1(n7227), .Y(n7240) );
  CLKBUFX3 U7281 ( .A(n9511), .Y(n8370) );
  OR2X1 U7282 ( .A(n2585), .B(n9338), .Y(n7241) );
  OR2X1 U7283 ( .A(n2584), .B(n9338), .Y(n7242) );
  OR2X1 U7284 ( .A(n2583), .B(n9338), .Y(n7243) );
  OR2X1 U7285 ( .A(n2582), .B(n9338), .Y(n7244) );
  NAND2X1 U7286 ( .A(n9373), .B(n9341), .Y(n7245) );
  OR2X1 U7287 ( .A(n2582), .B(n9339), .Y(n7246) );
  NAND2X1 U7288 ( .A(n9391), .B(n9362), .Y(n7247) );
  NAND2X1 U7289 ( .A(n2211), .B(n9342), .Y(n7248) );
  NAND2XL U7290 ( .A(n9459), .B(n1459), .Y(n1421) );
  DLY4X1 U7291 ( .A(n7251), .Y(n7250) );
  DLY4X1 U7292 ( .A(\buff[61][7] ), .Y(n7251) );
  BUFX2 U7293 ( .A(n7250), .Y(n7249) );
  DLY4X1 U7294 ( .A(n7254), .Y(n7253) );
  DLY4X1 U7295 ( .A(n2594), .Y(n7254) );
  BUFX2 U7296 ( .A(n7253), .Y(n7252) );
  OAI2BB1XL U7297 ( .A0N(\buff[63][0] ), .A1N(n9458), .B0(n99), .Y(n2594) );
  BUFX2 U7298 ( .A(n7256), .Y(n7255) );
  DLY4X4 U7299 ( .A(n7257), .Y(n7256) );
  DLY4X4 U7300 ( .A(n2595), .Y(n7257) );
  OAI2BB1XL U7301 ( .A0N(\buff[63][1] ), .A1N(n9458), .B0(n103), .Y(n2595) );
  BUFX2 U7302 ( .A(n7259), .Y(n7258) );
  DLY4X4 U7303 ( .A(n7260), .Y(n7259) );
  DLY4X4 U7304 ( .A(n2596), .Y(n7260) );
  OAI2BB1XL U7305 ( .A0N(\buff[63][2] ), .A1N(n9458), .B0(n106), .Y(n2596) );
  BUFX2 U7306 ( .A(n7262), .Y(n7261) );
  DLY4X4 U7307 ( .A(n7263), .Y(n7262) );
  DLY4X4 U7308 ( .A(n2597), .Y(n7263) );
  OAI2BB1XL U7309 ( .A0N(\buff[63][3] ), .A1N(n9458), .B0(n109), .Y(n2597) );
  DLY4X1 U7310 ( .A(\buff[63][4] ), .Y(n7265) );
  BUFX2 U7311 ( .A(n7265), .Y(n7264) );
  DLY4X4 U7312 ( .A(n2598), .Y(n7266) );
  OAI2BB1XL U7313 ( .A0N(n7264), .A1N(n9458), .B0(n112), .Y(n2598) );
  BUFX2 U7314 ( .A(n2599), .Y(n7267) );
  DLY4X4 U7315 ( .A(n7269), .Y(n7268) );
  OAI2BB1XL U7316 ( .A0N(n7268), .A1N(n9458), .B0(n115), .Y(n2599) );
  DLY4X1 U7317 ( .A(n7272), .Y(n7271) );
  DLY4X1 U7318 ( .A(\buff[56][6] ), .Y(n7272) );
  BUFX2 U7319 ( .A(n7271), .Y(n7270) );
  DLY4X1 U7320 ( .A(n7275), .Y(n7274) );
  DLY4X1 U7321 ( .A(\buff[56][7] ), .Y(n7275) );
  BUFX2 U7322 ( .A(n7274), .Y(n7273) );
  DLY4X1 U7323 ( .A(n7278), .Y(n7277) );
  DLY4X1 U7324 ( .A(n2602), .Y(n7278) );
  BUFX2 U7325 ( .A(n7277), .Y(n7276) );
  DLY4X1 U7326 ( .A(n7281), .Y(n7280) );
  DLY4X1 U7327 ( .A(n2603), .Y(n7281) );
  BUFX2 U7328 ( .A(n7280), .Y(n7279) );
  DLY4X1 U7329 ( .A(n7284), .Y(n7283) );
  DLY4X1 U7330 ( .A(n2604), .Y(n7284) );
  BUFX2 U7331 ( .A(n7283), .Y(n7282) );
  DLY4X1 U7332 ( .A(n2605), .Y(n7287) );
  BUFX2 U7333 ( .A(n7286), .Y(n7285) );
  DLY4X4 U7334 ( .A(n7287), .Y(n7286) );
  DLY4X1 U7335 ( .A(n2606), .Y(n7290) );
  BUFX2 U7336 ( .A(n7290), .Y(n7288) );
  DLY4X4 U7337 ( .A(\buff[62][4] ), .Y(n7289) );
  DLY4X1 U7338 ( .A(n7293), .Y(n7292) );
  DLY4X1 U7339 ( .A(\buff[62][5] ), .Y(n7293) );
  BUFX2 U7340 ( .A(n7292), .Y(n7291) );
  DLY4X1 U7341 ( .A(n7296), .Y(n7295) );
  DLY4X1 U7342 ( .A(\buff[59][6] ), .Y(n7296) );
  BUFX2 U7343 ( .A(n7295), .Y(n7294) );
  OAI2BB2X2 U7344 ( .B0(n9454), .B1(n185), .A0N(n7298), .A1N(n9454), .Y(n2633)
         );
  BUFX2 U7345 ( .A(n2633), .Y(n7297) );
  DLY4X4 U7346 ( .A(n7299), .Y(n7298) );
  DLY4X1 U7347 ( .A(n7302), .Y(n7301) );
  DLY4X1 U7348 ( .A(n2610), .Y(n7302) );
  BUFX2 U7349 ( .A(n7301), .Y(n7300) );
  DLY4X1 U7350 ( .A(n7305), .Y(n7304) );
  DLY4X1 U7351 ( .A(n2611), .Y(n7305) );
  BUFX2 U7352 ( .A(n7304), .Y(n7303) );
  DLY4X1 U7353 ( .A(n7308), .Y(n7307) );
  DLY4X1 U7354 ( .A(n2612), .Y(n7308) );
  BUFX2 U7355 ( .A(n7307), .Y(n7306) );
  DLY4X1 U7356 ( .A(n2613), .Y(n7311) );
  BUFX2 U7357 ( .A(n7310), .Y(n7309) );
  DLY4X4 U7358 ( .A(n7311), .Y(n7310) );
  DLY4X1 U7359 ( .A(n2614), .Y(n7314) );
  BUFX2 U7360 ( .A(n7314), .Y(n7312) );
  DLY4X4 U7361 ( .A(\buff[61][4] ), .Y(n7313) );
  DLY4X1 U7362 ( .A(n7317), .Y(n7316) );
  DLY4X1 U7363 ( .A(\buff[61][5] ), .Y(n7317) );
  BUFX2 U7364 ( .A(n7316), .Y(n7315) );
  DLY4X1 U7365 ( .A(n7320), .Y(n7319) );
  DLY4X1 U7366 ( .A(\buff[62][6] ), .Y(n7320) );
  BUFX2 U7367 ( .A(n7319), .Y(n7318) );
  DLY4X1 U7368 ( .A(n7323), .Y(n7322) );
  DLY4X1 U7369 ( .A(\buff[62][7] ), .Y(n7323) );
  BUFX2 U7370 ( .A(n7322), .Y(n7321) );
  DLY4X1 U7371 ( .A(n7326), .Y(n7325) );
  DLY4X1 U7372 ( .A(n2618), .Y(n7326) );
  BUFX2 U7373 ( .A(n7325), .Y(n7324) );
  DLY4X1 U7374 ( .A(n7329), .Y(n7328) );
  DLY4X1 U7375 ( .A(n2619), .Y(n7329) );
  BUFX2 U7376 ( .A(n7328), .Y(n7327) );
  DLY4X1 U7377 ( .A(n7332), .Y(n7331) );
  DLY4X1 U7378 ( .A(n2620), .Y(n7332) );
  BUFX2 U7379 ( .A(n7331), .Y(n7330) );
  DLY4X1 U7380 ( .A(n2621), .Y(n7335) );
  BUFX2 U7381 ( .A(n7334), .Y(n7333) );
  DLY4X4 U7382 ( .A(n7335), .Y(n7334) );
  DLY4X1 U7383 ( .A(n2622), .Y(n7338) );
  BUFX2 U7384 ( .A(n7338), .Y(n7336) );
  DLY4X4 U7385 ( .A(\buff[60][4] ), .Y(n7337) );
  DLY4X1 U7386 ( .A(n7341), .Y(n7340) );
  DLY4X1 U7387 ( .A(\buff[60][5] ), .Y(n7341) );
  BUFX2 U7388 ( .A(n7340), .Y(n7339) );
  DLY4X1 U7389 ( .A(n7344), .Y(n7343) );
  DLY4X1 U7390 ( .A(\buff[57][6] ), .Y(n7344) );
  BUFX2 U7391 ( .A(n7343), .Y(n7342) );
  DLY4X1 U7392 ( .A(n7347), .Y(n7346) );
  DLY4X1 U7393 ( .A(\buff[57][7] ), .Y(n7347) );
  BUFX2 U7394 ( .A(n7346), .Y(n7345) );
  BUFX2 U7395 ( .A(n7349), .Y(n7348) );
  DLY4X4 U7396 ( .A(n7350), .Y(n7349) );
  DLY4X4 U7397 ( .A(n2626), .Y(n7350) );
  BUFX2 U7398 ( .A(n7352), .Y(n7351) );
  DLY4X4 U7399 ( .A(n7353), .Y(n7352) );
  DLY4X4 U7400 ( .A(n2627), .Y(n7353) );
  BUFX2 U7401 ( .A(n7355), .Y(n7354) );
  DLY4X4 U7402 ( .A(n7356), .Y(n7355) );
  DLY4X4 U7403 ( .A(n2628), .Y(n7356) );
  BUFX2 U7404 ( .A(n7358), .Y(n7357) );
  DLY4X4 U7405 ( .A(n7359), .Y(n7358) );
  DLY4X4 U7406 ( .A(n2629), .Y(n7359) );
  DLY4X1 U7407 ( .A(\buff[59][4] ), .Y(n7361) );
  BUFX2 U7408 ( .A(n7361), .Y(n7360) );
  BUFX2 U7409 ( .A(n2631), .Y(n7363) );
  OA22XL U7410 ( .A0(n159), .A1(n186), .B0(n187), .B1(n145), .Y(n175) );
  DLY4X4 U7411 ( .A(n7365), .Y(n7364) );
  DLY4X1 U7412 ( .A(n7367), .Y(n7366) );
  DLY4X1 U7413 ( .A(n1413), .Y(n7367) );
  NAND2XL U7414 ( .A(\buff[28][6] ), .B(n9693), .Y(n1413) );
  DLY4X1 U7415 ( .A(n7369), .Y(n7368) );
  DLY4X1 U7416 ( .A(n1417), .Y(n7369) );
  NAND2XL U7417 ( .A(\buff[28][7] ), .B(n9693), .Y(n1417) );
  DLY4X1 U7418 ( .A(n7372), .Y(n7371) );
  DLY4X1 U7419 ( .A(n2634), .Y(n7372) );
  BUFX2 U7420 ( .A(n7371), .Y(n7370) );
  DLY4X1 U7421 ( .A(n7375), .Y(n7374) );
  DLY4X1 U7422 ( .A(n2635), .Y(n7375) );
  BUFX2 U7423 ( .A(n7374), .Y(n7373) );
  DLY4X1 U7424 ( .A(n7378), .Y(n7377) );
  DLY4X1 U7425 ( .A(n2636), .Y(n7378) );
  BUFX2 U7426 ( .A(n7377), .Y(n7376) );
  DLY4X1 U7427 ( .A(n2637), .Y(n7381) );
  BUFX2 U7428 ( .A(n7380), .Y(n7379) );
  DLY4X4 U7429 ( .A(n7381), .Y(n7380) );
  DLY4X1 U7430 ( .A(n2638), .Y(n7384) );
  BUFX2 U7431 ( .A(n7384), .Y(n7382) );
  DLY4X4 U7432 ( .A(\buff[58][4] ), .Y(n7383) );
  DLY4X1 U7433 ( .A(n7387), .Y(n7386) );
  DLY4X1 U7434 ( .A(\buff[58][5] ), .Y(n7387) );
  BUFX2 U7435 ( .A(n7386), .Y(n7385) );
  DLY4X1 U7436 ( .A(n7390), .Y(n7389) );
  DLY4X1 U7437 ( .A(\buff[60][6] ), .Y(n7390) );
  BUFX2 U7438 ( .A(n7389), .Y(n7388) );
  DLY4X1 U7439 ( .A(n7393), .Y(n7392) );
  DLY4X1 U7440 ( .A(\buff[60][7] ), .Y(n7393) );
  BUFX2 U7441 ( .A(n7392), .Y(n7391) );
  DLY4X1 U7442 ( .A(n7396), .Y(n7395) );
  DLY4X1 U7443 ( .A(n2642), .Y(n7396) );
  BUFX2 U7444 ( .A(n7395), .Y(n7394) );
  DLY4X1 U7445 ( .A(n7399), .Y(n7398) );
  DLY4X1 U7446 ( .A(n2643), .Y(n7399) );
  BUFX2 U7447 ( .A(n7398), .Y(n7397) );
  DLY4X1 U7448 ( .A(n7402), .Y(n7401) );
  DLY4X1 U7449 ( .A(n2644), .Y(n7402) );
  BUFX2 U7450 ( .A(n7401), .Y(n7400) );
  DLY4X1 U7451 ( .A(n2645), .Y(n7405) );
  BUFX2 U7452 ( .A(n7404), .Y(n7403) );
  DLY4X4 U7453 ( .A(n7405), .Y(n7404) );
  DLY4X1 U7454 ( .A(n2646), .Y(n7408) );
  BUFX2 U7455 ( .A(n7408), .Y(n7406) );
  DLY4X4 U7456 ( .A(\buff[57][4] ), .Y(n7407) );
  DLY4X1 U7457 ( .A(n7411), .Y(n7410) );
  DLY4X1 U7458 ( .A(\buff[57][5] ), .Y(n7411) );
  BUFX2 U7459 ( .A(n7410), .Y(n7409) );
  DLY4X1 U7460 ( .A(n7414), .Y(n7413) );
  DLY4X1 U7461 ( .A(\buff[58][6] ), .Y(n7414) );
  BUFX2 U7462 ( .A(n7413), .Y(n7412) );
  DLY4X1 U7463 ( .A(n7417), .Y(n7416) );
  DLY4X1 U7464 ( .A(\buff[58][7] ), .Y(n7417) );
  BUFX2 U7465 ( .A(n7416), .Y(n7415) );
  DLY4X1 U7466 ( .A(n7420), .Y(n7419) );
  DLY4X1 U7467 ( .A(n2650), .Y(n7420) );
  BUFX2 U7468 ( .A(n7419), .Y(n7418) );
  DLY4X1 U7469 ( .A(n7423), .Y(n7422) );
  DLY4X1 U7470 ( .A(n2651), .Y(n7423) );
  BUFX2 U7471 ( .A(n7422), .Y(n7421) );
  DLY4X1 U7472 ( .A(n7426), .Y(n7425) );
  DLY4X1 U7473 ( .A(n2652), .Y(n7426) );
  BUFX2 U7474 ( .A(n7425), .Y(n7424) );
  DLY4X1 U7475 ( .A(n2653), .Y(n7429) );
  BUFX2 U7476 ( .A(n7428), .Y(n7427) );
  DLY4X4 U7477 ( .A(n7429), .Y(n7428) );
  DLY4X1 U7478 ( .A(n2654), .Y(n7432) );
  BUFX2 U7479 ( .A(n7432), .Y(n7430) );
  DLY4X4 U7480 ( .A(\buff[56][4] ), .Y(n7431) );
  DLY4X1 U7481 ( .A(n7435), .Y(n7434) );
  DLY4X1 U7482 ( .A(\buff[56][5] ), .Y(n7435) );
  BUFX2 U7483 ( .A(n7434), .Y(n7433) );
  DLY4X1 U7484 ( .A(n1614), .Y(n7436) );
  DLY4X4 U7485 ( .A(n2921), .Y(n7437) );
  OAI211XL U7486 ( .A0(n9393), .A1(n288), .B0(n1613), .C0(n7436), .Y(n2921) );
  NAND2XL U7487 ( .A(\buff[23][7] ), .B(n9393), .Y(n1614) );
  DLY4X4 U7488 ( .A(n7439), .Y(n7438) );
  DLY4X4 U7489 ( .A(n7441), .Y(n7440) );
  DLY4X1 U7490 ( .A(n7443), .Y(n7442) );
  DLY4X4 U7491 ( .A(n2660), .Y(n7443) );
  DLY4X1 U7492 ( .A(n7445), .Y(n7444) );
  DLY4X4 U7493 ( .A(n2661), .Y(n7445) );
  DLY4X4 U7494 ( .A(\buff[55][4] ), .Y(n7446) );
  DLY4X4 U7495 ( .A(n2662), .Y(n7447) );
  DLY4X4 U7496 ( .A(n7449), .Y(n7448) );
  DLY4X4 U7497 ( .A(\buff[55][5] ), .Y(n7449) );
  DLY4X1 U7498 ( .A(n7451), .Y(n7450) );
  DLY4X1 U7499 ( .A(n2526), .Y(n7451) );
  NAND2XL U7500 ( .A(\buff[0][6] ), .B(n9670), .Y(n2526) );
  DLY4X1 U7501 ( .A(n7453), .Y(n7452) );
  DLY4X1 U7502 ( .A(n2530), .Y(n7453) );
  NAND2XL U7503 ( .A(\buff[0][7] ), .B(n9670), .Y(n2530) );
  DLY4X1 U7504 ( .A(n2666), .Y(n7454) );
  DLY4X1 U7505 ( .A(n304), .Y(n7455) );
  NAND2XL U7506 ( .A(\buff[54][0] ), .B(n9709), .Y(n304) );
  DLY4X1 U7507 ( .A(n2667), .Y(n7456) );
  DLY4X1 U7508 ( .A(n315), .Y(n7457) );
  NAND2XL U7509 ( .A(\buff[54][1] ), .B(n9709), .Y(n315) );
  DLY4X1 U7510 ( .A(n2668), .Y(n7458) );
  DLY4X1 U7511 ( .A(n323), .Y(n7459) );
  NAND2XL U7512 ( .A(\buff[54][2] ), .B(n9709), .Y(n323) );
  DLY4X1 U7513 ( .A(n2669), .Y(n7460) );
  DLY4X1 U7514 ( .A(n331), .Y(n7461) );
  NAND2XL U7515 ( .A(\buff[54][3] ), .B(n9709), .Y(n331) );
  DLY4X1 U7516 ( .A(n2670), .Y(n7462) );
  DLY4X1 U7517 ( .A(n339), .Y(n7463) );
  NAND2XL U7518 ( .A(\buff[54][4] ), .B(n9709), .Y(n339) );
  DLY4X1 U7519 ( .A(n2671), .Y(n7464) );
  DLY4X1 U7520 ( .A(n347), .Y(n7465) );
  NAND2XL U7521 ( .A(\buff[54][5] ), .B(n9709), .Y(n347) );
  DLY4X1 U7522 ( .A(n7467), .Y(n7466) );
  DLY4X1 U7523 ( .A(n2485), .Y(n7467) );
  NAND2XL U7524 ( .A(\buff[1][6] ), .B(n9677), .Y(n2485) );
  DLY4X1 U7525 ( .A(n7469), .Y(n7468) );
  DLY4X1 U7526 ( .A(n2489), .Y(n7469) );
  NAND2XL U7527 ( .A(\buff[1][7] ), .B(n9677), .Y(n2489) );
  DLY4X1 U7528 ( .A(n2674), .Y(n7470) );
  DLY4X1 U7529 ( .A(n379), .Y(n7471) );
  NAND2XL U7530 ( .A(\buff[53][0] ), .B(n9703), .Y(n379) );
  DLY4X1 U7531 ( .A(n2675), .Y(n7472) );
  DLY4X1 U7532 ( .A(n386), .Y(n7473) );
  NAND2XL U7533 ( .A(\buff[53][1] ), .B(n9703), .Y(n386) );
  BUFX12 U7534 ( .A(n2584), .Y(n7474) );
  OAI221X4 U7535 ( .A0(n389), .A1(n377), .B0(n9703), .B1(n9644), .C0(n7475), 
        .Y(n2676) );
  DLY4X1 U7536 ( .A(n7476), .Y(n7475) );
  DLY4X1 U7537 ( .A(n390), .Y(n7476) );
  NAND2XL U7538 ( .A(\buff[53][2] ), .B(n9703), .Y(n390) );
  DLY4X1 U7539 ( .A(n2677), .Y(n7477) );
  OAI221X2 U7540 ( .A0(n393), .A1(n377), .B0(n9703), .B1(n9641), .C0(n7478), 
        .Y(n2677) );
  DLY4X1 U7541 ( .A(n394), .Y(n7478) );
  NAND2XL U7542 ( .A(\buff[53][3] ), .B(n9703), .Y(n394) );
  DLY4X1 U7543 ( .A(n2678), .Y(n7479) );
  OAI221X2 U7544 ( .A0(n397), .A1(n377), .B0(n9703), .B1(n267), .C0(n7480), 
        .Y(n2678) );
  DLY4X1 U7545 ( .A(n398), .Y(n7480) );
  NAND2XL U7546 ( .A(\buff[53][4] ), .B(n9703), .Y(n398) );
  DLY4X1 U7547 ( .A(n2679), .Y(n7481) );
  OAI221X2 U7548 ( .A0(n401), .A1(n377), .B0(n9703), .B1(n9629), .C0(n7482), 
        .Y(n2679) );
  DLY4X1 U7549 ( .A(n402), .Y(n7482) );
  NAND2XL U7550 ( .A(\buff[53][5] ), .B(n9703), .Y(n402) );
  OAI221X4 U7551 ( .A0(n2282), .A1(n2255), .B0(n9704), .B1(n9625), .C0(n7483), 
        .Y(n3056) );
  DLY4X1 U7552 ( .A(n7484), .Y(n7483) );
  DLY4X1 U7553 ( .A(n2283), .Y(n7484) );
  NAND2XL U7554 ( .A(\buff[6][6] ), .B(n9704), .Y(n2283) );
  OAI221X4 U7555 ( .A0(n2286), .A1(n2255), .B0(n9704), .B1(n9618), .C0(n7485), 
        .Y(n3057) );
  DLY4X1 U7556 ( .A(n7486), .Y(n7485) );
  DLY4X1 U7557 ( .A(n2287), .Y(n7486) );
  NAND2XL U7558 ( .A(\buff[6][7] ), .B(n9704), .Y(n2287) );
  DLY4X1 U7559 ( .A(n2682), .Y(n7487) );
  DLY4X1 U7560 ( .A(n419), .Y(n7488) );
  NAND2XL U7561 ( .A(\buff[52][0] ), .B(n9696), .Y(n419) );
  OAI221X4 U7562 ( .A0(n425), .A1(n417), .B0(n9696), .B1(n9649), .C0(n7489), 
        .Y(n2683) );
  DLY4X1 U7563 ( .A(n7490), .Y(n7489) );
  DLY4X1 U7564 ( .A(n426), .Y(n7490) );
  NAND2XL U7565 ( .A(\buff[52][1] ), .B(n9696), .Y(n426) );
  OAI221X4 U7566 ( .A0(n429), .A1(n417), .B0(n9696), .B1(n9644), .C0(n7491), 
        .Y(n2684) );
  DLY4X1 U7567 ( .A(n7492), .Y(n7491) );
  DLY4X1 U7568 ( .A(n430), .Y(n7492) );
  NAND2XL U7569 ( .A(\buff[52][2] ), .B(n9696), .Y(n430) );
  DLY4X1 U7570 ( .A(n2685), .Y(n7493) );
  OAI221X2 U7571 ( .A0(n433), .A1(n417), .B0(n9696), .B1(n9641), .C0(n7494), 
        .Y(n2685) );
  DLY4X1 U7572 ( .A(n434), .Y(n7494) );
  NAND2XL U7573 ( .A(\buff[52][3] ), .B(n9696), .Y(n434) );
  DLY4X1 U7574 ( .A(n2686), .Y(n7495) );
  OAI221X2 U7575 ( .A0(n437), .A1(n417), .B0(n9696), .B1(n9635), .C0(n7496), 
        .Y(n2686) );
  DLY4X1 U7576 ( .A(n438), .Y(n7496) );
  NAND2XL U7577 ( .A(\buff[52][4] ), .B(n9696), .Y(n438) );
  DLY4X1 U7578 ( .A(n2687), .Y(n7497) );
  OAI221X2 U7579 ( .A0(n441), .A1(n417), .B0(n9696), .B1(n9629), .C0(n7498), 
        .Y(n2687) );
  DLY4X1 U7580 ( .A(n442), .Y(n7498) );
  NAND2XL U7581 ( .A(\buff[52][5] ), .B(n9696), .Y(n442) );
  DLY4X1 U7582 ( .A(n7500), .Y(n7499) );
  DLY4X1 U7583 ( .A(n7502), .Y(n7501) );
  DLY4X1 U7584 ( .A(n3108), .Y(n7502) );
  DLY4X1 U7585 ( .A(n2690), .Y(n7503) );
  OAI221XL U7586 ( .A0(n456), .A1(n457), .B0(n9689), .B1(n9656), .C0(n7504), 
        .Y(n2690) );
  DLY4X1 U7587 ( .A(n459), .Y(n7504) );
  NAND2XL U7588 ( .A(\buff[51][0] ), .B(n9689), .Y(n459) );
  DLY4X1 U7589 ( .A(n2691), .Y(n7505) );
  OAI221X2 U7590 ( .A0(n465), .A1(n457), .B0(n9689), .B1(n9650), .C0(n7506), 
        .Y(n2691) );
  DLY4X1 U7591 ( .A(n466), .Y(n7506) );
  NAND2XL U7592 ( .A(\buff[51][1] ), .B(n9689), .Y(n466) );
  DLY4X1 U7593 ( .A(n2692), .Y(n7507) );
  OAI221X2 U7594 ( .A0(n469), .A1(n457), .B0(n9689), .B1(n9643), .C0(n7508), 
        .Y(n2692) );
  DLY4X1 U7595 ( .A(n470), .Y(n7508) );
  NAND2XL U7596 ( .A(\buff[51][2] ), .B(n9689), .Y(n470) );
  DLY4X1 U7597 ( .A(n2693), .Y(n7509) );
  OAI221X2 U7598 ( .A0(n473), .A1(n457), .B0(n9689), .B1(n9640), .C0(n7510), 
        .Y(n2693) );
  DLY4X1 U7599 ( .A(n474), .Y(n7510) );
  NAND2XL U7600 ( .A(\buff[51][3] ), .B(n9689), .Y(n474) );
  DLY4X1 U7601 ( .A(n7512), .Y(n7511) );
  DLY4X1 U7602 ( .A(n2326), .Y(n7512) );
  NAND2XL U7603 ( .A(\buff[5][6] ), .B(n9697), .Y(n2326) );
  DLY4X1 U7604 ( .A(n7514), .Y(n7513) );
  DLY4X1 U7605 ( .A(n2330), .Y(n7514) );
  NAND2XL U7606 ( .A(\buff[5][7] ), .B(n9697), .Y(n2330) );
  DLY4X1 U7607 ( .A(n2698), .Y(n7515) );
  DLY4X1 U7608 ( .A(n499), .Y(n7516) );
  NAND2XL U7609 ( .A(\buff[50][0] ), .B(n9716), .Y(n499) );
  OAI221X4 U7610 ( .A0(n505), .A1(n7521), .B0(n9716), .B1(n9648), .C0(n7517), 
        .Y(n2699) );
  DLY4X1 U7611 ( .A(n7518), .Y(n7517) );
  NAND2X1 U7612 ( .A(\buff[50][1] ), .B(n9716), .Y(n506) );
  DLY4X1 U7613 ( .A(n506), .Y(n7518) );
  OAI221X4 U7614 ( .A0(n509), .A1(n7521), .B0(n9716), .B1(n9642), .C0(n7519), 
        .Y(n2700) );
  DLY4X1 U7615 ( .A(n7520), .Y(n7519) );
  NAND2X1 U7616 ( .A(\buff[50][2] ), .B(n9716), .Y(n510) );
  DLY4X1 U7617 ( .A(n510), .Y(n7520) );
  NAND2X1 U7618 ( .A(n9663), .B(n531), .Y(n497) );
  BUFX2 U7619 ( .A(n497), .Y(n7521) );
  OAI221X4 U7620 ( .A0(n513), .A1(n7521), .B0(n9716), .B1(n9639), .C0(n7522), 
        .Y(n2701) );
  DLY4X1 U7621 ( .A(n7523), .Y(n7522) );
  DLY4X1 U7622 ( .A(n514), .Y(n7523) );
  NAND2XL U7623 ( .A(\buff[50][3] ), .B(n9716), .Y(n514) );
  DLY4X1 U7624 ( .A(n2702), .Y(n7524) );
  OAI221X2 U7625 ( .A0(n517), .A1(n497), .B0(n9716), .B1(n9635), .C0(n7525), 
        .Y(n2702) );
  DLY4X1 U7626 ( .A(n518), .Y(n7525) );
  NAND2XL U7627 ( .A(\buff[50][4] ), .B(n9716), .Y(n518) );
  DLY4X1 U7628 ( .A(n2703), .Y(n7526) );
  OAI221X2 U7629 ( .A0(n521), .A1(n497), .B0(n9716), .B1(n9627), .C0(n7527), 
        .Y(n2703) );
  DLY4X1 U7630 ( .A(n522), .Y(n7527) );
  NAND2XL U7631 ( .A(\buff[50][5] ), .B(n9716), .Y(n522) );
  DLY4X4 U7632 ( .A(n7529), .Y(n7528) );
  DLY4X4 U7633 ( .A(\buff[55][6] ), .Y(n7529) );
  DLY4X4 U7634 ( .A(n7531), .Y(n7530) );
  DLY4X4 U7635 ( .A(\buff[55][7] ), .Y(n7531) );
  DLY4X1 U7636 ( .A(n2706), .Y(n7532) );
  DLY4X1 U7637 ( .A(n539), .Y(n7533) );
  NAND2XL U7638 ( .A(\buff[49][0] ), .B(n9683), .Y(n539) );
  DLY4X1 U7639 ( .A(n2707), .Y(n7534) );
  DLY4X1 U7640 ( .A(n546), .Y(n7535) );
  NAND2XL U7641 ( .A(\buff[49][1] ), .B(n9683), .Y(n546) );
  DLY4X1 U7642 ( .A(n2708), .Y(n7536) );
  DLY4X1 U7643 ( .A(n550), .Y(n7537) );
  NAND2XL U7644 ( .A(\buff[49][2] ), .B(n9683), .Y(n550) );
  BUFX2 U7645 ( .A(n537), .Y(n7538) );
  OAI221X4 U7646 ( .A0(n553), .A1(n7538), .B0(n9683), .B1(n9639), .C0(n7539), 
        .Y(n2709) );
  DLY4X1 U7647 ( .A(n7540), .Y(n7539) );
  DLY4X1 U7648 ( .A(n554), .Y(n7540) );
  NAND2XL U7649 ( .A(\buff[49][3] ), .B(n9683), .Y(n554) );
  DLY4X1 U7650 ( .A(n2710), .Y(n7541) );
  OAI221X2 U7651 ( .A0(n557), .A1(n537), .B0(n9683), .B1(n9635), .C0(n7542), 
        .Y(n2710) );
  DLY4X1 U7652 ( .A(n558), .Y(n7542) );
  NAND2XL U7653 ( .A(\buff[49][4] ), .B(n9683), .Y(n558) );
  DLY4X1 U7654 ( .A(n2711), .Y(n7543) );
  OAI221X2 U7655 ( .A0(n561), .A1(n537), .B0(n9683), .B1(n9627), .C0(n7544), 
        .Y(n2711) );
  DLY4X1 U7656 ( .A(n562), .Y(n7544) );
  NAND2XL U7657 ( .A(\buff[49][5] ), .B(n9683), .Y(n562) );
  DLY4X1 U7658 ( .A(n2445), .Y(n7545) );
  DLY4X4 U7659 ( .A(n3088), .Y(n7546) );
  OAI211XL U7660 ( .A0(n9625), .A1(n9360), .B0(n2444), .C0(n7545), .Y(n3088)
         );
  NAND2XL U7661 ( .A(\buff[2][6] ), .B(n9360), .Y(n2445) );
  DLY4X1 U7662 ( .A(\buff[2][7] ), .Y(n7547) );
  OAI211XL U7663 ( .A0(n9618), .A1(n9360), .B0(n2448), .C0(n2449), .Y(n3089)
         );
  NAND2XL U7664 ( .A(n7547), .B(n9360), .Y(n2449) );
  DLY4X1 U7665 ( .A(n2714), .Y(n7549) );
  DLY4X1 U7666 ( .A(n579), .Y(n7550) );
  NAND2XL U7667 ( .A(\buff[48][0] ), .B(n9676), .Y(n579) );
  OAI221X4 U7668 ( .A0(n585), .A1(n577), .B0(n9676), .B1(n9650), .C0(n7551), 
        .Y(n2715) );
  DLY4X1 U7669 ( .A(n7552), .Y(n7551) );
  DLY4X1 U7670 ( .A(n586), .Y(n7552) );
  NAND2XL U7671 ( .A(\buff[48][1] ), .B(n9676), .Y(n586) );
  OAI221X4 U7672 ( .A0(n589), .A1(n577), .B0(n9676), .B1(n9644), .C0(n7553), 
        .Y(n2716) );
  DLY4X1 U7673 ( .A(n7554), .Y(n7553) );
  DLY4X1 U7674 ( .A(n590), .Y(n7554) );
  NAND2XL U7675 ( .A(\buff[48][2] ), .B(n9676), .Y(n590) );
  DLY4X1 U7676 ( .A(n2717), .Y(n7555) );
  OAI221X2 U7677 ( .A0(n593), .A1(n577), .B0(n9676), .B1(n9641), .C0(n7556), 
        .Y(n2717) );
  DLY4X1 U7678 ( .A(n594), .Y(n7556) );
  NAND2XL U7679 ( .A(\buff[48][3] ), .B(n9676), .Y(n594) );
  DLY4X1 U7680 ( .A(n2718), .Y(n7557) );
  OAI221X2 U7681 ( .A0(n597), .A1(n577), .B0(n9676), .B1(n267), .C0(n7558), 
        .Y(n2718) );
  DLY4X1 U7682 ( .A(n598), .Y(n7558) );
  NAND2XL U7683 ( .A(\buff[48][4] ), .B(n9676), .Y(n598) );
  DLY4X1 U7684 ( .A(n2719), .Y(n7559) );
  OAI221X2 U7685 ( .A0(n601), .A1(n577), .B0(n9676), .B1(n9629), .C0(n7560), 
        .Y(n2719) );
  DLY4X1 U7686 ( .A(n602), .Y(n7560) );
  NAND2XL U7687 ( .A(\buff[48][5] ), .B(n9676), .Y(n602) );
  DLY4X1 U7688 ( .A(n3078), .Y(n7561) );
  OAI221XL U7689 ( .A0(n2397), .A1(n2376), .B0(n9684), .B1(n9634), .C0(n7562), 
        .Y(n3078) );
  DLY4X1 U7690 ( .A(n2398), .Y(n7562) );
  NAND2XL U7691 ( .A(\buff[3][4] ), .B(n9684), .Y(n2398) );
  DLY4X1 U7692 ( .A(n3079), .Y(n7563) );
  OAI221X2 U7693 ( .A0(n2401), .A1(n2376), .B0(n9684), .B1(n9628), .C0(n7564), 
        .Y(n3079) );
  DLY4X1 U7694 ( .A(n2402), .Y(n7564) );
  NAND2XL U7695 ( .A(\buff[3][5] ), .B(n9684), .Y(n2402) );
  DLY4X1 U7696 ( .A(n3080), .Y(n7565) );
  OAI221X2 U7697 ( .A0(n2405), .A1(n2376), .B0(n9684), .B1(n281), .C0(n7566), 
        .Y(n3080) );
  DLY4X1 U7698 ( .A(n2406), .Y(n7566) );
  NAND2XL U7699 ( .A(\buff[3][6] ), .B(n9684), .Y(n2406) );
  DLY4X1 U7700 ( .A(n3081), .Y(n7567) );
  OAI221X2 U7701 ( .A0(n2409), .A1(n2376), .B0(n9684), .B1(n9619), .C0(n7568), 
        .Y(n3081) );
  DLY4X1 U7702 ( .A(n2410), .Y(n7568) );
  NAND2XL U7703 ( .A(\buff[3][7] ), .B(n9684), .Y(n2410) );
  DLY4X1 U7704 ( .A(n7570), .Y(n7569) );
  OAI211XL U7705 ( .A0(n9423), .A1(n9655), .B0(n619), .C0(n620), .Y(n2722) );
  NAND2XL U7706 ( .A(\buff[47][0] ), .B(n9423), .Y(n620) );
  DLY4X1 U7707 ( .A(\buff[47][1] ), .Y(n7571) );
  OAI211XL U7708 ( .A0(n9423), .A1(n9650), .B0(n628), .C0(n629), .Y(n2723) );
  NAND2XL U7709 ( .A(n7571), .B(n9423), .Y(n629) );
  DLY4X1 U7710 ( .A(\buff[47][2] ), .Y(n7573) );
  OAI211XL U7711 ( .A0(n9423), .A1(n9644), .B0(n633), .C0(n634), .Y(n2724) );
  NAND2XL U7712 ( .A(n7573), .B(n9423), .Y(n634) );
  DLY4X1 U7713 ( .A(\buff[47][3] ), .Y(n7575) );
  OAI211XL U7714 ( .A0(n9423), .A1(n9641), .B0(n638), .C0(n639), .Y(n2725) );
  NAND2XL U7715 ( .A(n7575), .B(n9423), .Y(n639) );
  DLY4X1 U7716 ( .A(n2672), .Y(n7577) );
  OAI221X2 U7717 ( .A0(n354), .A1(n302), .B0(n9709), .B1(n9625), .C0(n7578), 
        .Y(n2672) );
  DLY4X1 U7718 ( .A(n355), .Y(n7578) );
  NAND2XL U7719 ( .A(\buff[54][6] ), .B(n9709), .Y(n355) );
  DLY4X1 U7720 ( .A(n2673), .Y(n7579) );
  OAI221X2 U7721 ( .A0(n362), .A1(n302), .B0(n9709), .B1(n9618), .C0(n7580), 
        .Y(n2673) );
  DLY4X1 U7722 ( .A(n363), .Y(n7580) );
  NAND2XL U7723 ( .A(\buff[54][7] ), .B(n9709), .Y(n363) );
  DLY4X1 U7724 ( .A(n2730), .Y(n7581) );
  DLY4X1 U7725 ( .A(n671), .Y(n7582) );
  NAND2XL U7726 ( .A(\buff[46][0] ), .B(n9708), .Y(n671) );
  DLY4X1 U7727 ( .A(n2731), .Y(n7583) );
  DLY4X1 U7728 ( .A(n678), .Y(n7584) );
  NAND2XL U7729 ( .A(\buff[46][1] ), .B(n9708), .Y(n678) );
  DLY4X1 U7730 ( .A(n2732), .Y(n7585) );
  DLY4X1 U7731 ( .A(n682), .Y(n7586) );
  NAND2XL U7732 ( .A(\buff[46][2] ), .B(n9708), .Y(n682) );
  DLY4X1 U7733 ( .A(n2733), .Y(n7587) );
  DLY4X1 U7734 ( .A(n686), .Y(n7588) );
  NAND2XL U7735 ( .A(\buff[46][3] ), .B(n9708), .Y(n686) );
  DLY4X1 U7736 ( .A(n2734), .Y(n7589) );
  DLY4X1 U7737 ( .A(n690), .Y(n7590) );
  NAND2XL U7738 ( .A(\buff[46][4] ), .B(n9708), .Y(n690) );
  DLY4X1 U7739 ( .A(n2735), .Y(n7591) );
  DLY4X1 U7740 ( .A(n694), .Y(n7592) );
  NAND2XL U7741 ( .A(\buff[46][5] ), .B(n9708), .Y(n694) );
  DLY4X4 U7742 ( .A(n2680), .Y(n7593) );
  OAI221X2 U7743 ( .A0(n405), .A1(n377), .B0(n9703), .B1(n9626), .C0(n7594), 
        .Y(n2680) );
  DLY4X1 U7744 ( .A(n406), .Y(n7594) );
  NAND2XL U7745 ( .A(\buff[53][6] ), .B(n9703), .Y(n406) );
  DLY4X1 U7746 ( .A(n2681), .Y(n7595) );
  OAI221X2 U7747 ( .A0(n409), .A1(n377), .B0(n9703), .B1(n9620), .C0(n7596), 
        .Y(n2681) );
  DLY4X1 U7748 ( .A(n410), .Y(n7596) );
  NAND2XL U7749 ( .A(\buff[53][7] ), .B(n9703), .Y(n410) );
  DLY4X1 U7750 ( .A(n2738), .Y(n7597) );
  DLY4X1 U7751 ( .A(n712), .Y(n7598) );
  NAND2XL U7752 ( .A(\buff[45][0] ), .B(n9702), .Y(n712) );
  DLY4X1 U7753 ( .A(n2739), .Y(n7599) );
  DLY4X1 U7754 ( .A(n719), .Y(n7600) );
  NAND2XL U7755 ( .A(\buff[45][1] ), .B(n9702), .Y(n719) );
  DLY4X1 U7756 ( .A(n2740), .Y(n7601) );
  DLY4X1 U7757 ( .A(n723), .Y(n7602) );
  NAND2XL U7758 ( .A(\buff[45][2] ), .B(n9702), .Y(n723) );
  DLY4X1 U7759 ( .A(n2741), .Y(n7603) );
  DLY4X1 U7760 ( .A(n727), .Y(n7604) );
  NAND2XL U7761 ( .A(\buff[45][3] ), .B(n9702), .Y(n727) );
  DLY4X1 U7762 ( .A(n2742), .Y(n7605) );
  DLY4X1 U7763 ( .A(n731), .Y(n7606) );
  NAND2XL U7764 ( .A(\buff[45][4] ), .B(n9702), .Y(n731) );
  DLY4X1 U7765 ( .A(n2743), .Y(n7607) );
  DLY4X1 U7766 ( .A(n735), .Y(n7608) );
  NAND2XL U7767 ( .A(\buff[45][5] ), .B(n9702), .Y(n735) );
  DLY4X4 U7768 ( .A(n2688), .Y(n7609) );
  OAI221X2 U7769 ( .A0(n445), .A1(n417), .B0(n9696), .B1(n9624), .C0(n7610), 
        .Y(n2688) );
  DLY4X1 U7770 ( .A(n446), .Y(n7610) );
  NAND2XL U7771 ( .A(\buff[52][6] ), .B(n9696), .Y(n446) );
  DLY4X1 U7772 ( .A(n2689), .Y(n7611) );
  OAI221X2 U7773 ( .A0(n449), .A1(n417), .B0(n9696), .B1(n9619), .C0(n7612), 
        .Y(n2689) );
  DLY4X1 U7774 ( .A(n450), .Y(n7612) );
  NAND2XL U7775 ( .A(\buff[52][7] ), .B(n9696), .Y(n450) );
  DLY4X1 U7776 ( .A(n2746), .Y(n7613) );
  DLY4X1 U7777 ( .A(n751), .Y(n7614) );
  NAND2XL U7778 ( .A(\buff[44][0] ), .B(n9695), .Y(n751) );
  DLY4X1 U7779 ( .A(n2747), .Y(n7615) );
  DLY4X1 U7780 ( .A(n758), .Y(n7616) );
  NAND2XL U7781 ( .A(\buff[44][1] ), .B(n9695), .Y(n758) );
  DLY4X1 U7782 ( .A(n2748), .Y(n7617) );
  DLY4X1 U7783 ( .A(n762), .Y(n7618) );
  NAND2XL U7784 ( .A(\buff[44][2] ), .B(n9695), .Y(n762) );
  DLY4X1 U7785 ( .A(n2749), .Y(n7619) );
  DLY4X1 U7786 ( .A(n766), .Y(n7620) );
  NAND2XL U7787 ( .A(\buff[44][3] ), .B(n9695), .Y(n766) );
  DLY4X1 U7788 ( .A(n2750), .Y(n7621) );
  DLY4X1 U7789 ( .A(n770), .Y(n7622) );
  NAND2XL U7790 ( .A(\buff[44][4] ), .B(n9695), .Y(n770) );
  DLY4X1 U7791 ( .A(n2751), .Y(n7623) );
  DLY4X1 U7792 ( .A(n774), .Y(n7624) );
  NAND2XL U7793 ( .A(\buff[44][5] ), .B(n9695), .Y(n774) );
  DLY4X1 U7794 ( .A(n2694), .Y(n7625) );
  OAI221X2 U7795 ( .A0(n477), .A1(n457), .B0(n9689), .B1(n9635), .C0(n7626), 
        .Y(n2694) );
  DLY4X1 U7796 ( .A(n478), .Y(n7626) );
  NAND2XL U7797 ( .A(\buff[51][4] ), .B(n9689), .Y(n478) );
  DLY4X1 U7798 ( .A(n2695), .Y(n7627) );
  OAI221X2 U7799 ( .A0(n481), .A1(n457), .B0(n9689), .B1(n9627), .C0(n7628), 
        .Y(n2695) );
  DLY4X1 U7800 ( .A(n482), .Y(n7628) );
  NAND2XL U7801 ( .A(\buff[51][5] ), .B(n9689), .Y(n482) );
  DLY4X1 U7802 ( .A(n2696), .Y(n7629) );
  OAI221X2 U7803 ( .A0(n485), .A1(n457), .B0(n9689), .B1(n281), .C0(n7630), 
        .Y(n2696) );
  DLY4X1 U7804 ( .A(n486), .Y(n7630) );
  NAND2XL U7805 ( .A(\buff[51][6] ), .B(n9689), .Y(n486) );
  DLY4X1 U7806 ( .A(n2697), .Y(n7631) );
  OAI221X2 U7807 ( .A0(n489), .A1(n457), .B0(n9689), .B1(n9619), .C0(n7632), 
        .Y(n2697) );
  DLY4X1 U7808 ( .A(n490), .Y(n7632) );
  NAND2XL U7809 ( .A(\buff[51][7] ), .B(n9689), .Y(n490) );
  DLY4X1 U7810 ( .A(n2754), .Y(n7633) );
  OAI221XL U7811 ( .A0(n787), .A1(n788), .B0(n9688), .B1(n9656), .C0(n7634), 
        .Y(n2754) );
  DLY4X1 U7812 ( .A(n790), .Y(n7634) );
  NAND2XL U7813 ( .A(\buff[43][0] ), .B(n9688), .Y(n790) );
  DLY4X1 U7814 ( .A(n2755), .Y(n7635) );
  OAI221X2 U7815 ( .A0(n796), .A1(n788), .B0(n9688), .B1(n9650), .C0(n7636), 
        .Y(n2755) );
  DLY4X1 U7816 ( .A(n797), .Y(n7636) );
  NAND2XL U7817 ( .A(\buff[43][1] ), .B(n9688), .Y(n797) );
  DLY4X1 U7818 ( .A(n2756), .Y(n7637) );
  OAI221X2 U7819 ( .A0(n800), .A1(n788), .B0(n9688), .B1(n9644), .C0(n7638), 
        .Y(n2756) );
  DLY4X1 U7820 ( .A(n801), .Y(n7638) );
  NAND2XL U7821 ( .A(\buff[43][2] ), .B(n9688), .Y(n801) );
  DLY4X1 U7822 ( .A(n2757), .Y(n7639) );
  OAI221X2 U7823 ( .A0(n804), .A1(n788), .B0(n9688), .B1(n9641), .C0(n7640), 
        .Y(n2757) );
  DLY4X1 U7824 ( .A(n805), .Y(n7640) );
  NAND2XL U7825 ( .A(\buff[43][3] ), .B(n9688), .Y(n805) );
  DLY4X4 U7826 ( .A(n2704), .Y(n7641) );
  OAI221X2 U7827 ( .A0(n525), .A1(n497), .B0(n9716), .B1(n9624), .C0(n7642), 
        .Y(n2704) );
  DLY4X1 U7828 ( .A(n526), .Y(n7642) );
  NAND2XL U7829 ( .A(\buff[50][6] ), .B(n9716), .Y(n526) );
  DLY4X1 U7830 ( .A(n2705), .Y(n7643) );
  OAI221X2 U7831 ( .A0(n529), .A1(n497), .B0(n9716), .B1(n9619), .C0(n7644), 
        .Y(n2705) );
  DLY4X1 U7832 ( .A(n530), .Y(n7644) );
  NAND2XL U7833 ( .A(\buff[50][7] ), .B(n9716), .Y(n530) );
  DLY4X1 U7834 ( .A(n2762), .Y(n7645) );
  DLY4X1 U7835 ( .A(n829), .Y(n7646) );
  NAND2XL U7836 ( .A(\buff[42][0] ), .B(n9715), .Y(n829) );
  OAI221X4 U7837 ( .A0(n835), .A1(n827), .B0(n9715), .B1(n9650), .C0(n7647), 
        .Y(n2763) );
  DLY4X1 U7838 ( .A(n7648), .Y(n7647) );
  DLY4X1 U7839 ( .A(n836), .Y(n7648) );
  NAND2XL U7840 ( .A(\buff[42][1] ), .B(n9715), .Y(n836) );
  OAI221X4 U7841 ( .A0(n839), .A1(n827), .B0(n9715), .B1(n9644), .C0(n7649), 
        .Y(n2764) );
  DLY4X1 U7842 ( .A(n7650), .Y(n7649) );
  DLY4X1 U7843 ( .A(n840), .Y(n7650) );
  NAND2XL U7844 ( .A(\buff[42][2] ), .B(n9715), .Y(n840) );
  OAI221X4 U7845 ( .A0(n843), .A1(n827), .B0(n9715), .B1(n9641), .C0(n7651), 
        .Y(n2765) );
  DLY4X1 U7846 ( .A(n7652), .Y(n7651) );
  DLY4X1 U7847 ( .A(n844), .Y(n7652) );
  NAND2XL U7848 ( .A(\buff[42][3] ), .B(n9715), .Y(n844) );
  OAI221X4 U7849 ( .A0(n847), .A1(n827), .B0(n9715), .B1(n9635), .C0(n7653), 
        .Y(n2766) );
  DLY4X1 U7850 ( .A(n7654), .Y(n7653) );
  DLY4X1 U7851 ( .A(n848), .Y(n7654) );
  NAND2XL U7852 ( .A(\buff[42][4] ), .B(n9715), .Y(n848) );
  OAI221X4 U7853 ( .A0(n851), .A1(n827), .B0(n9715), .B1(n9629), .C0(n7655), 
        .Y(n2767) );
  DLY4X1 U7854 ( .A(n7656), .Y(n7655) );
  DLY4X1 U7855 ( .A(n852), .Y(n7656) );
  NAND2XL U7856 ( .A(\buff[42][5] ), .B(n9715), .Y(n852) );
  DLY4X1 U7857 ( .A(n2712), .Y(n7657) );
  OAI221X2 U7858 ( .A0(n565), .A1(n537), .B0(n9683), .B1(n281), .C0(n7658), 
        .Y(n2712) );
  DLY4X1 U7859 ( .A(n566), .Y(n7658) );
  NAND2XL U7860 ( .A(\buff[49][6] ), .B(n9683), .Y(n566) );
  DLY4X1 U7861 ( .A(n2713), .Y(n7659) );
  OAI221X2 U7862 ( .A0(n569), .A1(n537), .B0(n9683), .B1(n9618), .C0(n7660), 
        .Y(n2713) );
  DLY4X1 U7863 ( .A(n570), .Y(n7660) );
  NAND2XL U7864 ( .A(\buff[49][7] ), .B(n9683), .Y(n570) );
  DLY4X1 U7865 ( .A(n2770), .Y(n7661) );
  DLY4X1 U7866 ( .A(n868), .Y(n7662) );
  NAND2XL U7867 ( .A(\buff[41][0] ), .B(n9682), .Y(n868) );
  DLY4X1 U7868 ( .A(n2771), .Y(n7663) );
  DLY4X1 U7869 ( .A(n875), .Y(n7664) );
  NAND2XL U7870 ( .A(\buff[41][1] ), .B(n9682), .Y(n875) );
  DLY4X1 U7871 ( .A(n2772), .Y(n7665) );
  DLY4X1 U7872 ( .A(n879), .Y(n7666) );
  NAND2XL U7873 ( .A(\buff[41][2] ), .B(n9682), .Y(n879) );
  DLY4X1 U7874 ( .A(n2773), .Y(n7667) );
  DLY4X1 U7875 ( .A(n883), .Y(n7668) );
  NAND2XL U7876 ( .A(\buff[41][3] ), .B(n9682), .Y(n883) );
  DLY4X1 U7877 ( .A(n2774), .Y(n7669) );
  DLY4X1 U7878 ( .A(n887), .Y(n7670) );
  NAND2XL U7879 ( .A(\buff[41][4] ), .B(n9682), .Y(n887) );
  DLY4X1 U7880 ( .A(n2775), .Y(n7671) );
  DLY4X1 U7881 ( .A(n891), .Y(n7672) );
  NAND2XL U7882 ( .A(\buff[41][5] ), .B(n9682), .Y(n891) );
  DLY4X4 U7883 ( .A(n2720), .Y(n7673) );
  OAI221X2 U7884 ( .A0(n605), .A1(n577), .B0(n9676), .B1(n9626), .C0(n7674), 
        .Y(n2720) );
  DLY4X1 U7885 ( .A(n606), .Y(n7674) );
  NAND2XL U7886 ( .A(\buff[48][6] ), .B(n9676), .Y(n606) );
  DLY4X1 U7887 ( .A(n2721), .Y(n7675) );
  OAI221X2 U7888 ( .A0(n609), .A1(n577), .B0(n9676), .B1(n9620), .C0(n7676), 
        .Y(n2721) );
  DLY4X1 U7889 ( .A(n610), .Y(n7676) );
  NAND2XL U7890 ( .A(\buff[48][7] ), .B(n9676), .Y(n610) );
  DLY4X1 U7891 ( .A(n2778), .Y(n7677) );
  DLY4X1 U7892 ( .A(n907), .Y(n7678) );
  NAND2XL U7893 ( .A(\buff[40][0] ), .B(n9675), .Y(n907) );
  DLY4X1 U7894 ( .A(n2779), .Y(n7679) );
  DLY4X1 U7895 ( .A(n914), .Y(n7680) );
  NAND2XL U7896 ( .A(\buff[40][1] ), .B(n9675), .Y(n914) );
  DLY4X1 U7897 ( .A(n2780), .Y(n7681) );
  DLY4X1 U7898 ( .A(n918), .Y(n7682) );
  NAND2XL U7899 ( .A(\buff[40][2] ), .B(n9675), .Y(n918) );
  DLY4X1 U7900 ( .A(n2781), .Y(n7683) );
  DLY4X1 U7901 ( .A(n922), .Y(n7684) );
  NAND2XL U7902 ( .A(\buff[40][3] ), .B(n9675), .Y(n922) );
  DLY4X1 U7903 ( .A(n2782), .Y(n7685) );
  DLY4X1 U7904 ( .A(n926), .Y(n7686) );
  NAND2XL U7905 ( .A(\buff[40][4] ), .B(n9675), .Y(n926) );
  DLY4X1 U7906 ( .A(n2783), .Y(n7687) );
  DLY4X1 U7907 ( .A(n930), .Y(n7688) );
  NAND2XL U7908 ( .A(\buff[40][5] ), .B(n9675), .Y(n930) );
  DLY4X1 U7909 ( .A(\buff[47][4] ), .Y(n7689) );
  OAI211XL U7910 ( .A0(n9423), .A1(n9635), .B0(n643), .C0(n644), .Y(n2726) );
  NAND2XL U7911 ( .A(n7689), .B(n9423), .Y(n644) );
  DLY4X1 U7912 ( .A(\buff[47][5] ), .Y(n7691) );
  OAI211XL U7913 ( .A0(n9423), .A1(n9628), .B0(n648), .C0(n649), .Y(n2727) );
  NAND2XL U7914 ( .A(n7691), .B(n9423), .Y(n649) );
  DLY3X1 U7915 ( .A(n2728), .Y(n7693) );
  OAI211XL U7916 ( .A0(n9423), .A1(n9625), .B0(n653), .C0(n7694), .Y(n2728) );
  DLY4X1 U7917 ( .A(n654), .Y(n7694) );
  NAND2XL U7918 ( .A(\buff[47][6] ), .B(n9423), .Y(n654) );
  DLY4X1 U7919 ( .A(n659), .Y(n7695) );
  DLY4X4 U7920 ( .A(n2729), .Y(n7696) );
  OAI211XL U7921 ( .A0(n9423), .A1(n288), .B0(n658), .C0(n7695), .Y(n2729) );
  NAND2XL U7922 ( .A(\buff[47][7] ), .B(n9423), .Y(n659) );
  DLY4X1 U7923 ( .A(n7698), .Y(n7697) );
  OAI211XL U7924 ( .A0(n9654), .A1(n9413), .B0(n944), .C0(n945), .Y(n2786) );
  NAND2XL U7925 ( .A(\buff[39][0] ), .B(n9413), .Y(n945) );
  DLY4X1 U7926 ( .A(\buff[39][1] ), .Y(n7699) );
  OAI211XL U7927 ( .A0(n9649), .A1(n9413), .B0(n952), .C0(n953), .Y(n2787) );
  NAND2XL U7928 ( .A(n7699), .B(n9413), .Y(n953) );
  DLY4X1 U7929 ( .A(\buff[39][2] ), .Y(n7701) );
  OAI211XL U7930 ( .A0(n9643), .A1(n9413), .B0(n956), .C0(n957), .Y(n2788) );
  NAND2XL U7931 ( .A(n7701), .B(n9413), .Y(n957) );
  DLY4X1 U7932 ( .A(\buff[39][3] ), .Y(n7703) );
  OAI211XL U7933 ( .A0(n9640), .A1(n9413), .B0(n960), .C0(n961), .Y(n2789) );
  NAND2XL U7934 ( .A(n7703), .B(n9413), .Y(n961) );
  DLY4X1 U7935 ( .A(n7706), .Y(n7705) );
  DLY4X1 U7936 ( .A(n698), .Y(n7706) );
  NAND2XL U7937 ( .A(\buff[46][6] ), .B(n9708), .Y(n698) );
  DLY4X1 U7938 ( .A(n7708), .Y(n7707) );
  DLY4X1 U7939 ( .A(n702), .Y(n7708) );
  NAND2XL U7940 ( .A(\buff[46][7] ), .B(n9708), .Y(n702) );
  DLY4X1 U7941 ( .A(n2794), .Y(n7709) );
  DLY4X1 U7942 ( .A(n991), .Y(n7710) );
  NAND2XL U7943 ( .A(\buff[38][0] ), .B(n9707), .Y(n991) );
  DLY4X1 U7944 ( .A(n2795), .Y(n7711) );
  DLY4X1 U7945 ( .A(n998), .Y(n7712) );
  NAND2XL U7946 ( .A(\buff[38][1] ), .B(n9707), .Y(n998) );
  DLY4X1 U7947 ( .A(n2796), .Y(n7713) );
  DLY4X1 U7948 ( .A(n1002), .Y(n7714) );
  NAND2XL U7949 ( .A(\buff[38][2] ), .B(n9707), .Y(n1002) );
  DLY4X1 U7950 ( .A(n2797), .Y(n7715) );
  DLY4X1 U7951 ( .A(n1006), .Y(n7716) );
  NAND2XL U7952 ( .A(\buff[38][3] ), .B(n9707), .Y(n1006) );
  DLY4X1 U7953 ( .A(n2798), .Y(n7717) );
  DLY4X1 U7954 ( .A(n1010), .Y(n7718) );
  NAND2XL U7955 ( .A(\buff[38][4] ), .B(n9707), .Y(n1010) );
  DLY4X1 U7956 ( .A(n2799), .Y(n7719) );
  DLY4X1 U7957 ( .A(n1014), .Y(n7720) );
  NAND2XL U7958 ( .A(\buff[38][5] ), .B(n9707), .Y(n1014) );
  DLY4X1 U7959 ( .A(n7722), .Y(n7721) );
  DLY4X1 U7960 ( .A(n739), .Y(n7722) );
  NAND2XL U7961 ( .A(\buff[45][6] ), .B(n9702), .Y(n739) );
  DLY4X1 U7962 ( .A(n7724), .Y(n7723) );
  DLY4X1 U7963 ( .A(n743), .Y(n7724) );
  NAND2XL U7964 ( .A(\buff[45][7] ), .B(n9702), .Y(n743) );
  DLY4X1 U7965 ( .A(n2802), .Y(n7725) );
  DLY4X1 U7966 ( .A(n1032), .Y(n7726) );
  NAND2XL U7967 ( .A(\buff[37][0] ), .B(n9701), .Y(n1032) );
  DLY4X1 U7968 ( .A(n2803), .Y(n7727) );
  DLY4X1 U7969 ( .A(n1039), .Y(n7728) );
  NAND2XL U7970 ( .A(\buff[37][1] ), .B(n9701), .Y(n1039) );
  DLY4X1 U7971 ( .A(n2804), .Y(n7729) );
  DLY4X1 U7972 ( .A(n1043), .Y(n7730) );
  NAND2XL U7973 ( .A(\buff[37][2] ), .B(n9701), .Y(n1043) );
  DLY4X1 U7974 ( .A(n2805), .Y(n7731) );
  DLY4X1 U7975 ( .A(n1047), .Y(n7732) );
  NAND2XL U7976 ( .A(\buff[37][3] ), .B(n9701), .Y(n1047) );
  DLY4X1 U7977 ( .A(n2806), .Y(n7733) );
  DLY4X1 U7978 ( .A(n1051), .Y(n7734) );
  NAND2XL U7979 ( .A(\buff[37][4] ), .B(n9701), .Y(n1051) );
  DLY4X1 U7980 ( .A(n2807), .Y(n7735) );
  DLY4X1 U7981 ( .A(n1055), .Y(n7736) );
  NAND2XL U7982 ( .A(\buff[37][5] ), .B(n9701), .Y(n1055) );
  DLY4X1 U7983 ( .A(n7738), .Y(n7737) );
  DLY4X1 U7984 ( .A(n778), .Y(n7738) );
  NAND2XL U7985 ( .A(\buff[44][6] ), .B(n9695), .Y(n778) );
  DLY4X1 U7986 ( .A(n7740), .Y(n7739) );
  DLY4X1 U7987 ( .A(n782), .Y(n7740) );
  NAND2XL U7988 ( .A(\buff[44][7] ), .B(n9695), .Y(n782) );
  DLY4X1 U7989 ( .A(n2810), .Y(n7741) );
  DLY4X1 U7990 ( .A(n1071), .Y(n7742) );
  NAND2XL U7991 ( .A(\buff[36][0] ), .B(n9694), .Y(n1071) );
  DLY4X1 U7992 ( .A(n2811), .Y(n7743) );
  DLY4X1 U7993 ( .A(n1078), .Y(n7744) );
  NAND2XL U7994 ( .A(\buff[36][1] ), .B(n9694), .Y(n1078) );
  DLY4X1 U7995 ( .A(n2812), .Y(n7745) );
  DLY4X1 U7996 ( .A(n1082), .Y(n7746) );
  NAND2XL U7997 ( .A(\buff[36][2] ), .B(n9694), .Y(n1082) );
  DLY4X1 U7998 ( .A(n2813), .Y(n7747) );
  DLY4X1 U7999 ( .A(n1086), .Y(n7748) );
  NAND2XL U8000 ( .A(\buff[36][3] ), .B(n9694), .Y(n1086) );
  DLY4X1 U8001 ( .A(n2814), .Y(n7749) );
  DLY4X1 U8002 ( .A(n1090), .Y(n7750) );
  NAND2XL U8003 ( .A(\buff[36][4] ), .B(n9694), .Y(n1090) );
  DLY4X1 U8004 ( .A(n2815), .Y(n7751) );
  DLY4X1 U8005 ( .A(n1094), .Y(n7752) );
  NAND2XL U8006 ( .A(\buff[36][5] ), .B(n9694), .Y(n1094) );
  DLY4X1 U8007 ( .A(n2758), .Y(n7753) );
  OAI221X2 U8008 ( .A0(n808), .A1(n788), .B0(n9688), .B1(n267), .C0(n7754), 
        .Y(n2758) );
  DLY4X1 U8009 ( .A(n809), .Y(n7754) );
  NAND2XL U8010 ( .A(\buff[43][4] ), .B(n9688), .Y(n809) );
  DLY4X1 U8011 ( .A(n2759), .Y(n7755) );
  OAI221X2 U8012 ( .A0(n812), .A1(n788), .B0(n9688), .B1(n9629), .C0(n7756), 
        .Y(n2759) );
  DLY4X1 U8013 ( .A(n813), .Y(n7756) );
  NAND2XL U8014 ( .A(\buff[43][5] ), .B(n9688), .Y(n813) );
  DLY4X1 U8015 ( .A(n2760), .Y(n7757) );
  OAI221X2 U8016 ( .A0(n816), .A1(n788), .B0(n9688), .B1(n9626), .C0(n7758), 
        .Y(n2760) );
  DLY4X1 U8017 ( .A(n817), .Y(n7758) );
  NAND2XL U8018 ( .A(\buff[43][6] ), .B(n9688), .Y(n817) );
  DLY4X1 U8019 ( .A(n2761), .Y(n7759) );
  OAI221X2 U8020 ( .A0(n820), .A1(n788), .B0(n9688), .B1(n9620), .C0(n7760), 
        .Y(n2761) );
  DLY4X1 U8021 ( .A(n821), .Y(n7760) );
  NAND2XL U8022 ( .A(\buff[43][7] ), .B(n9688), .Y(n821) );
  DLY4X1 U8023 ( .A(n2818), .Y(n7761) );
  OAI221XL U8024 ( .A0(n1107), .A1(n1108), .B0(n9687), .B1(n9656), .C0(n7762), 
        .Y(n2818) );
  DLY4X1 U8025 ( .A(n1110), .Y(n7762) );
  NAND2XL U8026 ( .A(\buff[35][0] ), .B(n9687), .Y(n1110) );
  DLY4X1 U8027 ( .A(n2819), .Y(n7763) );
  OAI221X2 U8028 ( .A0(n1116), .A1(n1108), .B0(n9687), .B1(n9650), .C0(n7764), 
        .Y(n2819) );
  DLY4X1 U8029 ( .A(n1117), .Y(n7764) );
  NAND2XL U8030 ( .A(\buff[35][1] ), .B(n9687), .Y(n1117) );
  DLY4X1 U8031 ( .A(n2820), .Y(n7765) );
  OAI221X2 U8032 ( .A0(n1120), .A1(n1108), .B0(n9687), .B1(n9644), .C0(n7766), 
        .Y(n2820) );
  DLY4X1 U8033 ( .A(n1121), .Y(n7766) );
  NAND2XL U8034 ( .A(\buff[35][2] ), .B(n9687), .Y(n1121) );
  DLY4X1 U8035 ( .A(n2821), .Y(n7767) );
  OAI221X2 U8036 ( .A0(n1124), .A1(n1108), .B0(n9687), .B1(n9641), .C0(n7768), 
        .Y(n2821) );
  DLY4X1 U8037 ( .A(n1125), .Y(n7768) );
  NAND2XL U8038 ( .A(\buff[35][3] ), .B(n9687), .Y(n1125) );
  OAI221X4 U8039 ( .A0(n855), .A1(n827), .B0(n9715), .B1(n9626), .C0(n7769), 
        .Y(n2768) );
  DLY4X1 U8040 ( .A(n7770), .Y(n7769) );
  DLY4X1 U8041 ( .A(n856), .Y(n7770) );
  NAND2XL U8042 ( .A(\buff[42][6] ), .B(n9715), .Y(n856) );
  OAI221X4 U8043 ( .A0(n859), .A1(n827), .B0(n9715), .B1(n9620), .C0(n7771), 
        .Y(n2769) );
  DLY4X1 U8044 ( .A(n7772), .Y(n7771) );
  DLY4X1 U8045 ( .A(n860), .Y(n7772) );
  NAND2XL U8046 ( .A(\buff[42][7] ), .B(n9715), .Y(n860) );
  DLY4X1 U8047 ( .A(n2826), .Y(n7773) );
  DLY4X1 U8048 ( .A(n1149), .Y(n7774) );
  NAND2XL U8049 ( .A(\buff[34][0] ), .B(n9714), .Y(n1149) );
  DLY4X1 U8050 ( .A(n2827), .Y(n7775) );
  DLY4X1 U8051 ( .A(n1156), .Y(n7776) );
  NAND2XL U8052 ( .A(\buff[34][1] ), .B(n9714), .Y(n1156) );
  OAI221X4 U8053 ( .A0(n1159), .A1(n1147), .B0(n9714), .B1(n9644), .C0(n7777), 
        .Y(n2828) );
  DLY4X1 U8054 ( .A(n7778), .Y(n7777) );
  DLY4X1 U8055 ( .A(n1160), .Y(n7778) );
  NAND2XL U8056 ( .A(\buff[34][2] ), .B(n9714), .Y(n1160) );
  OAI221X4 U8057 ( .A0(n1163), .A1(n1147), .B0(n9714), .B1(n9641), .C0(n7779), 
        .Y(n2829) );
  DLY4X1 U8058 ( .A(n7780), .Y(n7779) );
  DLY4X1 U8059 ( .A(n1164), .Y(n7780) );
  NAND2XL U8060 ( .A(\buff[34][3] ), .B(n9714), .Y(n1164) );
  OAI221X4 U8061 ( .A0(n1167), .A1(n1147), .B0(n9714), .B1(n9635), .C0(n7781), 
        .Y(n2830) );
  DLY4X1 U8062 ( .A(n7782), .Y(n7781) );
  DLY4X1 U8063 ( .A(n1168), .Y(n7782) );
  NAND2XL U8064 ( .A(\buff[34][4] ), .B(n9714), .Y(n1168) );
  OAI221X4 U8065 ( .A0(n1171), .A1(n1147), .B0(n9714), .B1(n9629), .C0(n7783), 
        .Y(n2831) );
  DLY4X1 U8066 ( .A(n7784), .Y(n7783) );
  DLY4X1 U8067 ( .A(n1172), .Y(n7784) );
  NAND2XL U8068 ( .A(\buff[34][5] ), .B(n9714), .Y(n1172) );
  DLY4X1 U8069 ( .A(n7786), .Y(n7785) );
  DLY4X1 U8070 ( .A(n895), .Y(n7786) );
  NAND2XL U8071 ( .A(\buff[41][6] ), .B(n9682), .Y(n895) );
  DLY4X1 U8072 ( .A(n7788), .Y(n7787) );
  DLY4X1 U8073 ( .A(n899), .Y(n7788) );
  NAND2XL U8074 ( .A(\buff[41][7] ), .B(n9682), .Y(n899) );
  DLY4X1 U8075 ( .A(n2834), .Y(n7789) );
  DLY4X1 U8076 ( .A(n1188), .Y(n7790) );
  NAND2XL U8077 ( .A(\buff[33][0] ), .B(n9681), .Y(n1188) );
  DLY4X1 U8078 ( .A(n2835), .Y(n7791) );
  DLY4X1 U8079 ( .A(n1195), .Y(n7792) );
  NAND2XL U8080 ( .A(\buff[33][1] ), .B(n9681), .Y(n1195) );
  DLY4X1 U8081 ( .A(n2836), .Y(n7793) );
  DLY4X1 U8082 ( .A(n1199), .Y(n7794) );
  NAND2XL U8083 ( .A(\buff[33][2] ), .B(n9681), .Y(n1199) );
  DLY4X1 U8084 ( .A(n2837), .Y(n7795) );
  DLY4X1 U8085 ( .A(n1203), .Y(n7796) );
  NAND2XL U8086 ( .A(\buff[33][3] ), .B(n9681), .Y(n1203) );
  DLY4X1 U8087 ( .A(n2838), .Y(n7797) );
  DLY4X1 U8088 ( .A(n1207), .Y(n7798) );
  NAND2XL U8089 ( .A(\buff[33][4] ), .B(n9681), .Y(n1207) );
  DLY4X1 U8090 ( .A(n2839), .Y(n7799) );
  DLY4X1 U8091 ( .A(n1211), .Y(n7800) );
  NAND2XL U8092 ( .A(\buff[33][5] ), .B(n9681), .Y(n1211) );
  DLY4X1 U8093 ( .A(n7802), .Y(n7801) );
  DLY4X1 U8094 ( .A(n934), .Y(n7802) );
  NAND2XL U8095 ( .A(\buff[40][6] ), .B(n9675), .Y(n934) );
  DLY4X1 U8096 ( .A(n7804), .Y(n7803) );
  DLY4X1 U8097 ( .A(n938), .Y(n7804) );
  NAND2XL U8098 ( .A(\buff[40][7] ), .B(n9675), .Y(n938) );
  DLY4X1 U8099 ( .A(n2842), .Y(n7805) );
  DLY4X1 U8100 ( .A(n1227), .Y(n7806) );
  NAND2XL U8101 ( .A(\buff[32][0] ), .B(n9674), .Y(n1227) );
  BUFX2 U8102 ( .A(n1024), .Y(n7807) );
  OAI221X4 U8103 ( .A0(n1233), .A1(n1225), .B0(n9674), .B1(n9650), .C0(n7808), 
        .Y(n2843) );
  DLY4X1 U8104 ( .A(n7809), .Y(n7808) );
  NAND2X1 U8105 ( .A(\buff[32][1] ), .B(n9674), .Y(n1234) );
  DLY4X1 U8106 ( .A(n1234), .Y(n7809) );
  DLY4X1 U8107 ( .A(n2844), .Y(n7810) );
  OAI221X2 U8108 ( .A0(n1237), .A1(n1225), .B0(n9674), .B1(n9644), .C0(n7811), 
        .Y(n2844) );
  DLY4X1 U8109 ( .A(n1238), .Y(n7811) );
  NAND2XL U8110 ( .A(\buff[32][2] ), .B(n9674), .Y(n1238) );
  DLY4X1 U8111 ( .A(n2845), .Y(n7812) );
  OAI221X2 U8112 ( .A0(n1241), .A1(n1225), .B0(n9674), .B1(n9641), .C0(n7813), 
        .Y(n2845) );
  DLY4X1 U8113 ( .A(n1242), .Y(n7813) );
  NAND2XL U8114 ( .A(\buff[32][3] ), .B(n9674), .Y(n1242) );
  DLY4X1 U8115 ( .A(n2846), .Y(n7814) );
  OAI221X2 U8116 ( .A0(n1245), .A1(n1225), .B0(n9674), .B1(n9634), .C0(n7815), 
        .Y(n2846) );
  DLY4X1 U8117 ( .A(n1246), .Y(n7815) );
  NAND2XL U8118 ( .A(\buff[32][4] ), .B(n9674), .Y(n1246) );
  DLY4X1 U8119 ( .A(n2847), .Y(n7816) );
  OAI221X2 U8120 ( .A0(n1249), .A1(n1225), .B0(n9674), .B1(n9629), .C0(n7817), 
        .Y(n2847) );
  DLY4X1 U8121 ( .A(n1250), .Y(n7817) );
  NAND2XL U8122 ( .A(\buff[32][5] ), .B(n9674), .Y(n1250) );
  DLY4X1 U8123 ( .A(\buff[39][4] ), .Y(n7818) );
  OAI211XL U8124 ( .A0(n9633), .A1(n9413), .B0(n964), .C0(n965), .Y(n2790) );
  NAND2XL U8125 ( .A(n7818), .B(n9413), .Y(n965) );
  DLY4X1 U8126 ( .A(\buff[39][5] ), .Y(n7820) );
  OAI211XL U8127 ( .A0(n9627), .A1(n9413), .B0(n968), .C0(n969), .Y(n2791) );
  NAND2XL U8128 ( .A(n7820), .B(n9413), .Y(n969) );
  DLY3X1 U8129 ( .A(n2792), .Y(n7822) );
  OAI211X4 U8130 ( .A0(n9625), .A1(n9413), .B0(n972), .C0(n7823), .Y(n2792) );
  DLY4X1 U8131 ( .A(n973), .Y(n7823) );
  NAND2XL U8132 ( .A(\buff[39][6] ), .B(n9413), .Y(n973) );
  DLY4X1 U8133 ( .A(n977), .Y(n7824) );
  DLY4X4 U8134 ( .A(n2793), .Y(n7825) );
  OAI211XL U8135 ( .A0(n9618), .A1(n9413), .B0(n976), .C0(n7824), .Y(n2793) );
  NAND2XL U8136 ( .A(\buff[39][7] ), .B(n9413), .Y(n977) );
  DLY4X1 U8137 ( .A(n7827), .Y(n7826) );
  OAI211XL U8138 ( .A0(n9403), .A1(n9655), .B0(n1264), .C0(n1265), .Y(n2850)
         );
  NAND2XL U8139 ( .A(\buff[31][0] ), .B(n9403), .Y(n1265) );
  DLY4X1 U8140 ( .A(\buff[31][1] ), .Y(n7828) );
  OAI211XL U8141 ( .A0(n9403), .A1(n9650), .B0(n1272), .C0(n1273), .Y(n2851)
         );
  NAND2XL U8142 ( .A(n7828), .B(n9403), .Y(n1273) );
  DLY4X1 U8143 ( .A(\buff[31][2] ), .Y(n7830) );
  OAI211XL U8144 ( .A0(n9403), .A1(n9644), .B0(n1276), .C0(n1277), .Y(n2852)
         );
  NAND2XL U8145 ( .A(n7830), .B(n9403), .Y(n1277) );
  DLY4X1 U8146 ( .A(\buff[31][3] ), .Y(n7832) );
  OAI211XL U8147 ( .A0(n9403), .A1(n9641), .B0(n1280), .C0(n1281), .Y(n2853)
         );
  NAND2XL U8148 ( .A(n7832), .B(n9403), .Y(n1281) );
  DLY4X1 U8149 ( .A(n7835), .Y(n7834) );
  DLY4X1 U8150 ( .A(n1571), .Y(n7835) );
  NAND2XL U8151 ( .A(\buff[24][6] ), .B(n9673), .Y(n1571) );
  DLY4X1 U8152 ( .A(n7837), .Y(n7836) );
  DLY4X1 U8153 ( .A(n1575), .Y(n7837) );
  NAND2XL U8154 ( .A(\buff[24][7] ), .B(n9673), .Y(n1575) );
  DLY4X1 U8155 ( .A(n2858), .Y(n7838) );
  DLY4X1 U8156 ( .A(n1306), .Y(n7839) );
  NAND2XL U8157 ( .A(\buff[30][0] ), .B(n9706), .Y(n1306) );
  DLY4X1 U8158 ( .A(n2859), .Y(n7840) );
  DLY4X1 U8159 ( .A(n1313), .Y(n7841) );
  NAND2XL U8160 ( .A(\buff[30][1] ), .B(n9706), .Y(n1313) );
  DLY4X1 U8161 ( .A(n2860), .Y(n7842) );
  DLY4X1 U8162 ( .A(n1317), .Y(n7843) );
  NAND2XL U8163 ( .A(\buff[30][2] ), .B(n9706), .Y(n1317) );
  DLY4X1 U8164 ( .A(n2861), .Y(n7844) );
  DLY4X1 U8165 ( .A(n1321), .Y(n7845) );
  NAND2XL U8166 ( .A(\buff[30][3] ), .B(n9706), .Y(n1321) );
  DLY4X1 U8167 ( .A(n2862), .Y(n7846) );
  DLY4X1 U8168 ( .A(n1325), .Y(n7847) );
  NAND2XL U8169 ( .A(\buff[30][4] ), .B(n9706), .Y(n1325) );
  DLY4X1 U8170 ( .A(n2863), .Y(n7848) );
  DLY4X1 U8171 ( .A(n1329), .Y(n7849) );
  NAND2XL U8172 ( .A(\buff[30][5] ), .B(n9706), .Y(n1329) );
  DLY4X1 U8173 ( .A(n2808), .Y(n7850) );
  OAI221X2 U8174 ( .A0(n1058), .A1(n1030), .B0(n9701), .B1(n9626), .C0(n7851), 
        .Y(n2808) );
  DLY4X1 U8175 ( .A(n1059), .Y(n7851) );
  NAND2XL U8176 ( .A(\buff[37][6] ), .B(n9701), .Y(n1059) );
  DLY4X1 U8177 ( .A(n2809), .Y(n7852) );
  OAI221X2 U8178 ( .A0(n1062), .A1(n1030), .B0(n9701), .B1(n9620), .C0(n7853), 
        .Y(n2809) );
  DLY4X1 U8179 ( .A(n1063), .Y(n7853) );
  NAND2XL U8180 ( .A(\buff[37][7] ), .B(n9701), .Y(n1063) );
  DLY4X1 U8181 ( .A(n2866), .Y(n7854) );
  DLY4X1 U8182 ( .A(n1347), .Y(n7855) );
  NAND2XL U8183 ( .A(\buff[29][0] ), .B(n9700), .Y(n1347) );
  DLY4X1 U8184 ( .A(n2867), .Y(n7856) );
  DLY4X1 U8185 ( .A(n1354), .Y(n7857) );
  NAND2XL U8186 ( .A(\buff[29][1] ), .B(n9700), .Y(n1354) );
  DLY4X1 U8187 ( .A(n2868), .Y(n7858) );
  DLY4X1 U8188 ( .A(n1358), .Y(n7859) );
  NAND2XL U8189 ( .A(\buff[29][2] ), .B(n9700), .Y(n1358) );
  DLY4X1 U8190 ( .A(n2869), .Y(n7860) );
  DLY4X1 U8191 ( .A(n1362), .Y(n7861) );
  NAND2XL U8192 ( .A(\buff[29][3] ), .B(n9700), .Y(n1362) );
  DLY4X1 U8193 ( .A(n2870), .Y(n7862) );
  DLY4X1 U8194 ( .A(n1366), .Y(n7863) );
  NAND2XL U8195 ( .A(\buff[29][4] ), .B(n9700), .Y(n1366) );
  DLY4X1 U8196 ( .A(n2871), .Y(n7864) );
  DLY4X1 U8197 ( .A(n1370), .Y(n7865) );
  NAND2XL U8198 ( .A(\buff[29][5] ), .B(n9700), .Y(n1370) );
  DLY4X1 U8199 ( .A(n7867), .Y(n7866) );
  DLY4X1 U8200 ( .A(n1333), .Y(n7867) );
  NAND2XL U8201 ( .A(\buff[30][6] ), .B(n9706), .Y(n1333) );
  DLY4X1 U8202 ( .A(n7869), .Y(n7868) );
  DLY4X1 U8203 ( .A(n1337), .Y(n7869) );
  NAND2XL U8204 ( .A(\buff[30][7] ), .B(n9706), .Y(n1337) );
  DLY4X1 U8205 ( .A(n2874), .Y(n7870) );
  DLY4X1 U8206 ( .A(n1386), .Y(n7871) );
  NAND2XL U8207 ( .A(\buff[28][0] ), .B(n9693), .Y(n1386) );
  DLY4X1 U8208 ( .A(n2875), .Y(n7872) );
  DLY4X1 U8209 ( .A(n1393), .Y(n7873) );
  NAND2XL U8210 ( .A(\buff[28][1] ), .B(n9693), .Y(n1393) );
  DLY4X1 U8211 ( .A(n2876), .Y(n7874) );
  DLY4X1 U8212 ( .A(n1397), .Y(n7875) );
  NAND2XL U8213 ( .A(\buff[28][2] ), .B(n9693), .Y(n1397) );
  DLY4X1 U8214 ( .A(n2877), .Y(n7876) );
  DLY4X1 U8215 ( .A(n1401), .Y(n7877) );
  NAND2XL U8216 ( .A(\buff[28][3] ), .B(n9693), .Y(n1401) );
  DLY4X1 U8217 ( .A(n2878), .Y(n7878) );
  DLY4X1 U8218 ( .A(n1405), .Y(n7879) );
  NAND2XL U8219 ( .A(\buff[28][4] ), .B(n9693), .Y(n1405) );
  DLY4X1 U8220 ( .A(n2879), .Y(n7880) );
  DLY4X1 U8221 ( .A(n1409), .Y(n7881) );
  NAND2XL U8222 ( .A(\buff[28][5] ), .B(n9693), .Y(n1409) );
  DLY4X1 U8223 ( .A(n7883), .Y(n7882) );
  OAI211XL U8224 ( .A0(n9375), .A1(n9635), .B0(n2235), .C0(n2236), .Y(n3046)
         );
  NAND2XL U8225 ( .A(\buff[7][4] ), .B(n9375), .Y(n2236) );
  DLY4X1 U8226 ( .A(n2240), .Y(n7884) );
  DLY4X4 U8227 ( .A(n3047), .Y(n7885) );
  OAI211XL U8228 ( .A0(n9375), .A1(n9629), .B0(n2239), .C0(n7884), .Y(n3047)
         );
  NAND2XL U8229 ( .A(\buff[7][5] ), .B(n9375), .Y(n2240) );
  DLY4X1 U8230 ( .A(\buff[27][0] ), .Y(n7886) );
  OAI211XL U8231 ( .A0(n9654), .A1(n9397), .B0(n1422), .C0(n1423), .Y(n2882)
         );
  NAND2XL U8232 ( .A(n7886), .B(n9397), .Y(n1423) );
  DLY4X1 U8233 ( .A(\buff[27][1] ), .Y(n7888) );
  OAI211XL U8234 ( .A0(n9649), .A1(n9397), .B0(n1430), .C0(n1431), .Y(n2883)
         );
  NAND2XL U8235 ( .A(n7888), .B(n9397), .Y(n1431) );
  DLY4X1 U8236 ( .A(\buff[27][2] ), .Y(n7890) );
  OAI211XL U8237 ( .A0(n9643), .A1(n9397), .B0(n1434), .C0(n1435), .Y(n2884)
         );
  NAND2XL U8238 ( .A(n7890), .B(n9397), .Y(n1435) );
  DLY4X1 U8239 ( .A(\buff[27][3] ), .Y(n7892) );
  OAI211XL U8240 ( .A0(n9640), .A1(n9397), .B0(n1438), .C0(n1439), .Y(n2885)
         );
  NAND2XL U8241 ( .A(n7892), .B(n9397), .Y(n1439) );
  DLY4X1 U8242 ( .A(\buff[27][4] ), .Y(n7894) );
  OAI211XL U8243 ( .A0(n9633), .A1(n9397), .B0(n1442), .C0(n1443), .Y(n2886)
         );
  NAND2XL U8244 ( .A(n7894), .B(n9397), .Y(n1443) );
  DLY4X1 U8245 ( .A(\buff[27][5] ), .Y(n7896) );
  OAI211XL U8246 ( .A0(n9627), .A1(n9397), .B0(n1446), .C0(n1447), .Y(n2887)
         );
  NAND2XL U8247 ( .A(n7896), .B(n9397), .Y(n1447) );
  DLY4X1 U8248 ( .A(n7899), .Y(n7898) );
  DLY4X1 U8249 ( .A(n2366), .Y(n7899) );
  NAND2XL U8250 ( .A(\buff[4][6] ), .B(n9690), .Y(n2366) );
  DLY4X1 U8251 ( .A(n7901), .Y(n7900) );
  DLY4X1 U8252 ( .A(n2370), .Y(n7901) );
  NAND2XL U8253 ( .A(\buff[4][7] ), .B(n9690), .Y(n2370) );
  DLY4X1 U8254 ( .A(n2890), .Y(n7902) );
  DLY4X1 U8255 ( .A(n1466), .Y(n7903) );
  NAND2XL U8256 ( .A(\buff[26][0] ), .B(n9713), .Y(n1466) );
  OAI221X4 U8257 ( .A0(n1472), .A1(n1464), .B0(n9713), .B1(n9648), .C0(n7904), 
        .Y(n2891) );
  DLY4X1 U8258 ( .A(n7905), .Y(n7904) );
  DLY4X1 U8259 ( .A(n1473), .Y(n7905) );
  NAND2XL U8260 ( .A(\buff[26][1] ), .B(n9713), .Y(n1473) );
  OAI221X4 U8261 ( .A0(n1476), .A1(n1464), .B0(n9713), .B1(n9642), .C0(n7906), 
        .Y(n2892) );
  DLY4X1 U8262 ( .A(n7907), .Y(n7906) );
  DLY4X1 U8263 ( .A(n1477), .Y(n7907) );
  NAND2XL U8264 ( .A(\buff[26][2] ), .B(n9713), .Y(n1477) );
  OAI221X4 U8265 ( .A0(n1480), .A1(n1464), .B0(n9713), .B1(n9639), .C0(n7908), 
        .Y(n2893) );
  DLY4X1 U8266 ( .A(n7909), .Y(n7908) );
  DLY4X1 U8267 ( .A(n1481), .Y(n7909) );
  NAND2XL U8268 ( .A(\buff[26][3] ), .B(n9713), .Y(n1481) );
  OAI221X4 U8269 ( .A0(n1484), .A1(n1464), .B0(n9713), .B1(n9634), .C0(n7910), 
        .Y(n2894) );
  DLY4X1 U8270 ( .A(n7911), .Y(n7910) );
  DLY4X1 U8271 ( .A(n1485), .Y(n7911) );
  NAND2XL U8272 ( .A(\buff[26][4] ), .B(n9713), .Y(n1485) );
  OAI221X4 U8273 ( .A0(n1488), .A1(n1464), .B0(n9713), .B1(n9628), .C0(n7912), 
        .Y(n2895) );
  DLY4X1 U8274 ( .A(n7913), .Y(n7912) );
  DLY4X1 U8275 ( .A(n1489), .Y(n7913) );
  NAND2XL U8276 ( .A(\buff[26][5] ), .B(n9713), .Y(n1489) );
  DLY4X1 U8277 ( .A(n2840), .Y(n7914) );
  OAI221X2 U8278 ( .A0(n1214), .A1(n1186), .B0(n9681), .B1(n9626), .C0(n7915), 
        .Y(n2840) );
  DLY4X1 U8279 ( .A(n1215), .Y(n7915) );
  NAND2XL U8280 ( .A(\buff[33][6] ), .B(n9681), .Y(n1215) );
  DLY4X1 U8281 ( .A(n2841), .Y(n7916) );
  OAI221X2 U8282 ( .A0(n1218), .A1(n1186), .B0(n9681), .B1(n9620), .C0(n7917), 
        .Y(n2841) );
  DLY4X1 U8283 ( .A(n1219), .Y(n7917) );
  NAND2XL U8284 ( .A(\buff[33][7] ), .B(n9681), .Y(n1219) );
  DLY4X1 U8285 ( .A(n2898), .Y(n7918) );
  DLY4X1 U8286 ( .A(n1505), .Y(n7919) );
  NAND2XL U8287 ( .A(\buff[25][0] ), .B(n9680), .Y(n1505) );
  DLY4X1 U8288 ( .A(n2899), .Y(n7920) );
  DLY4X1 U8289 ( .A(n1512), .Y(n7921) );
  NAND2XL U8290 ( .A(\buff[25][1] ), .B(n9680), .Y(n1512) );
  DLY4X1 U8291 ( .A(n2900), .Y(n7922) );
  DLY4X1 U8292 ( .A(n1516), .Y(n7923) );
  NAND2XL U8293 ( .A(\buff[25][2] ), .B(n9680), .Y(n1516) );
  DLY4X1 U8294 ( .A(n2901), .Y(n7924) );
  DLY4X1 U8295 ( .A(n1520), .Y(n7925) );
  NAND2XL U8296 ( .A(\buff[25][3] ), .B(n9680), .Y(n1520) );
  DLY4X1 U8297 ( .A(n2902), .Y(n7926) );
  DLY4X1 U8298 ( .A(n1524), .Y(n7927) );
  NAND2XL U8299 ( .A(\buff[25][4] ), .B(n9680), .Y(n1524) );
  DLY4X1 U8300 ( .A(n2903), .Y(n7928) );
  DLY4X1 U8301 ( .A(n1528), .Y(n7929) );
  NAND2XL U8302 ( .A(\buff[25][5] ), .B(n9680), .Y(n1528) );
  OAI221X4 U8303 ( .A0(n1492), .A1(n1464), .B0(n9713), .B1(n9624), .C0(n7930), 
        .Y(n2896) );
  DLY4X1 U8304 ( .A(n7931), .Y(n7930) );
  DLY4X1 U8305 ( .A(n1493), .Y(n7931) );
  NAND2XL U8306 ( .A(\buff[26][6] ), .B(n9713), .Y(n1493) );
  OAI221X4 U8307 ( .A0(n1496), .A1(n1464), .B0(n9713), .B1(n9619), .C0(n7932), 
        .Y(n2897) );
  DLY4X1 U8308 ( .A(n7933), .Y(n7932) );
  DLY4X1 U8309 ( .A(n1497), .Y(n7933) );
  NAND2XL U8310 ( .A(\buff[26][7] ), .B(n9713), .Y(n1497) );
  DLY4X1 U8311 ( .A(n2906), .Y(n7934) );
  DLY4X1 U8312 ( .A(n1544), .Y(n7935) );
  NAND2XL U8313 ( .A(\buff[24][0] ), .B(n9673), .Y(n1544) );
  DLY4X1 U8314 ( .A(n2907), .Y(n7936) );
  DLY4X1 U8315 ( .A(n1551), .Y(n7937) );
  NAND2XL U8316 ( .A(\buff[24][1] ), .B(n9673), .Y(n1551) );
  DLY4X1 U8317 ( .A(n2908), .Y(n7938) );
  DLY4X1 U8318 ( .A(n1555), .Y(n7939) );
  NAND2XL U8319 ( .A(\buff[24][2] ), .B(n9673), .Y(n1555) );
  DLY4X1 U8320 ( .A(n2909), .Y(n7940) );
  DLY4X1 U8321 ( .A(n1559), .Y(n7941) );
  NAND2XL U8322 ( .A(\buff[24][3] ), .B(n9673), .Y(n1559) );
  DLY4X1 U8323 ( .A(n2910), .Y(n7942) );
  DLY4X1 U8324 ( .A(n1563), .Y(n7943) );
  NAND2XL U8325 ( .A(\buff[24][4] ), .B(n9673), .Y(n1563) );
  DLY4X1 U8326 ( .A(n2911), .Y(n7944) );
  DLY4X1 U8327 ( .A(n1567), .Y(n7945) );
  NAND2XL U8328 ( .A(\buff[24][5] ), .B(n9673), .Y(n1567) );
  DLY4X1 U8329 ( .A(\buff[27][6] ), .Y(n7946) );
  OAI211X4 U8330 ( .A0(n9625), .A1(n9397), .B0(n1450), .C0(n7947), .Y(n2888)
         );
  DLY4X1 U8331 ( .A(n1451), .Y(n7947) );
  NAND2XL U8332 ( .A(n7946), .B(n9397), .Y(n1451) );
  DLY4X1 U8333 ( .A(\buff[27][7] ), .Y(n7948) );
  OAI211XL U8334 ( .A0(n9618), .A1(n9397), .B0(n1454), .C0(n1455), .Y(n2889)
         );
  NAND2XL U8335 ( .A(n7948), .B(n9397), .Y(n1455) );
  DLY4X1 U8336 ( .A(n7951), .Y(n7950) );
  OAI211XL U8337 ( .A0(n9393), .A1(n9655), .B0(n1581), .C0(n1582), .Y(n2914)
         );
  NAND2XL U8338 ( .A(\buff[23][0] ), .B(n9393), .Y(n1582) );
  DLY4X1 U8339 ( .A(n7953), .Y(n7952) );
  OAI211XL U8340 ( .A0(n9393), .A1(n9648), .B0(n1589), .C0(n1590), .Y(n2915)
         );
  NAND2XL U8341 ( .A(\buff[23][1] ), .B(n9393), .Y(n1590) );
  DLY4X1 U8342 ( .A(n7955), .Y(n7954) );
  OAI211XL U8343 ( .A0(n9393), .A1(n9642), .B0(n1593), .C0(n1594), .Y(n2916)
         );
  NAND2XL U8344 ( .A(\buff[23][2] ), .B(n9393), .Y(n1594) );
  DLY4X1 U8345 ( .A(n7957), .Y(n7956) );
  OAI211XL U8346 ( .A0(n9393), .A1(n9639), .B0(n1597), .C0(n1598), .Y(n2917)
         );
  NAND2XL U8347 ( .A(\buff[23][3] ), .B(n9393), .Y(n1598) );
  DLY4X1 U8348 ( .A(n7959), .Y(n7958) );
  OAI211XL U8349 ( .A0(n9393), .A1(n9635), .B0(n1601), .C0(n1602), .Y(n2918)
         );
  NAND2XL U8350 ( .A(\buff[23][4] ), .B(n9393), .Y(n1602) );
  DLY4X1 U8351 ( .A(n1606), .Y(n7960) );
  DLY4X4 U8352 ( .A(n2919), .Y(n7961) );
  OAI211XL U8353 ( .A0(n9393), .A1(n9628), .B0(n1605), .C0(n7960), .Y(n2919)
         );
  NAND2XL U8354 ( .A(\buff[23][5] ), .B(n9393), .Y(n1606) );
  DLY4X1 U8355 ( .A(n2800), .Y(n7962) );
  OAI221X2 U8356 ( .A0(n1017), .A1(n989), .B0(n9707), .B1(n9626), .C0(n7963), 
        .Y(n2800) );
  DLY4X1 U8357 ( .A(n1018), .Y(n7963) );
  NAND2XL U8358 ( .A(\buff[38][6] ), .B(n9707), .Y(n1018) );
  DLY4X1 U8359 ( .A(n2801), .Y(n7964) );
  OAI221X2 U8360 ( .A0(n1021), .A1(n989), .B0(n9707), .B1(n9620), .C0(n7965), 
        .Y(n2801) );
  DLY4X1 U8361 ( .A(n1022), .Y(n7965) );
  NAND2XL U8362 ( .A(\buff[38][7] ), .B(n9707), .Y(n1022) );
  DLY4X1 U8363 ( .A(n2922), .Y(n7966) );
  DLY4X1 U8364 ( .A(n1622), .Y(n7967) );
  NAND2XL U8365 ( .A(\buff[22][0] ), .B(n9705), .Y(n1622) );
  DLY4X1 U8366 ( .A(n2923), .Y(n7968) );
  DLY4X1 U8367 ( .A(n1628), .Y(n7969) );
  NAND2XL U8368 ( .A(\buff[22][1] ), .B(n9705), .Y(n1628) );
  DLY4X1 U8369 ( .A(n2924), .Y(n7970) );
  DLY4X1 U8370 ( .A(n1632), .Y(n7971) );
  NAND2XL U8371 ( .A(\buff[22][2] ), .B(n9705), .Y(n1632) );
  DLY4X1 U8372 ( .A(n2925), .Y(n7972) );
  DLY4X1 U8373 ( .A(n1636), .Y(n7973) );
  NAND2XL U8374 ( .A(\buff[22][3] ), .B(n9705), .Y(n1636) );
  DLY4X1 U8375 ( .A(n2926), .Y(n7974) );
  DLY4X1 U8376 ( .A(n1640), .Y(n7975) );
  NAND2XL U8377 ( .A(\buff[22][4] ), .B(n9705), .Y(n1640) );
  DLY4X1 U8378 ( .A(n2927), .Y(n7976) );
  DLY4X1 U8379 ( .A(n1644), .Y(n7977) );
  NAND2XL U8380 ( .A(\buff[22][5] ), .B(n9705), .Y(n1644) );
  DLY4X1 U8381 ( .A(n7979), .Y(n7978) );
  DLY4X1 U8382 ( .A(n1374), .Y(n7979) );
  NAND2XL U8383 ( .A(\buff[29][6] ), .B(n9700), .Y(n1374) );
  DLY4X1 U8384 ( .A(n7981), .Y(n7980) );
  DLY4X1 U8385 ( .A(n1378), .Y(n7981) );
  NAND2XL U8386 ( .A(\buff[29][7] ), .B(n9700), .Y(n1378) );
  DLY4X1 U8387 ( .A(n2930), .Y(n7982) );
  DLY4X1 U8388 ( .A(n1662), .Y(n7983) );
  NAND2XL U8389 ( .A(\buff[21][0] ), .B(n9699), .Y(n1662) );
  DLY4X1 U8390 ( .A(n2931), .Y(n7984) );
  DLY4X1 U8391 ( .A(n1669), .Y(n7985) );
  NAND2XL U8392 ( .A(\buff[21][1] ), .B(n9699), .Y(n1669) );
  DLY4X1 U8393 ( .A(n2932), .Y(n7986) );
  DLY4X1 U8394 ( .A(n1673), .Y(n7987) );
  NAND2XL U8395 ( .A(\buff[21][2] ), .B(n9699), .Y(n1673) );
  DLY4X1 U8396 ( .A(n2933), .Y(n7988) );
  DLY4X1 U8397 ( .A(n1677), .Y(n7989) );
  NAND2XL U8398 ( .A(\buff[21][3] ), .B(n9699), .Y(n1677) );
  DLY4X1 U8399 ( .A(n2934), .Y(n7990) );
  DLY4X1 U8400 ( .A(n1681), .Y(n7991) );
  NAND2XL U8401 ( .A(\buff[21][4] ), .B(n9699), .Y(n1681) );
  DLY4X1 U8402 ( .A(n2935), .Y(n7992) );
  DLY4X1 U8403 ( .A(n1685), .Y(n7993) );
  NAND2XL U8404 ( .A(\buff[21][5] ), .B(n9699), .Y(n1685) );
  DLY4X1 U8405 ( .A(n2816), .Y(n7994) );
  OAI221X2 U8406 ( .A0(n1097), .A1(n1069), .B0(n9694), .B1(n9626), .C0(n7995), 
        .Y(n2816) );
  DLY4X1 U8407 ( .A(n1098), .Y(n7995) );
  NAND2XL U8408 ( .A(\buff[36][6] ), .B(n9694), .Y(n1098) );
  DLY4X1 U8409 ( .A(n2817), .Y(n7996) );
  OAI221X2 U8410 ( .A0(n1101), .A1(n1069), .B0(n9694), .B1(n9620), .C0(n7997), 
        .Y(n2817) );
  DLY4X1 U8411 ( .A(n1102), .Y(n7997) );
  NAND2XL U8412 ( .A(\buff[36][7] ), .B(n9694), .Y(n1102) );
  DLY4X1 U8413 ( .A(n2938), .Y(n7998) );
  DLY4X1 U8414 ( .A(n1701), .Y(n7999) );
  NAND2XL U8415 ( .A(\buff[20][0] ), .B(n9692), .Y(n1701) );
  DLY4X1 U8416 ( .A(n2939), .Y(n8000) );
  DLY4X1 U8417 ( .A(n1708), .Y(n8001) );
  NAND2XL U8418 ( .A(\buff[20][1] ), .B(n9692), .Y(n1708) );
  DLY4X1 U8419 ( .A(n2940), .Y(n8002) );
  DLY4X1 U8420 ( .A(n1712), .Y(n8003) );
  NAND2XL U8421 ( .A(\buff[20][2] ), .B(n9692), .Y(n1712) );
  DLY4X1 U8422 ( .A(n2941), .Y(n8004) );
  DLY4X1 U8423 ( .A(n1716), .Y(n8005) );
  NAND2XL U8424 ( .A(\buff[20][3] ), .B(n9692), .Y(n1716) );
  DLY4X1 U8425 ( .A(n2942), .Y(n8006) );
  DLY4X1 U8426 ( .A(n1720), .Y(n8007) );
  NAND2XL U8427 ( .A(\buff[20][4] ), .B(n9692), .Y(n1720) );
  DLY4X1 U8428 ( .A(n2943), .Y(n8008) );
  DLY4X1 U8429 ( .A(n1724), .Y(n8009) );
  NAND2XL U8430 ( .A(\buff[20][5] ), .B(n9692), .Y(n1724) );
  DLY4X1 U8431 ( .A(n2822), .Y(n8010) );
  OAI221X2 U8432 ( .A0(n1128), .A1(n1108), .B0(n9687), .B1(n9635), .C0(n8011), 
        .Y(n2822) );
  DLY4X1 U8433 ( .A(n1129), .Y(n8011) );
  NAND2XL U8434 ( .A(\buff[35][4] ), .B(n9687), .Y(n1129) );
  DLY4X1 U8435 ( .A(n2823), .Y(n8012) );
  OAI221X2 U8436 ( .A0(n1132), .A1(n1108), .B0(n9687), .B1(n9629), .C0(n8013), 
        .Y(n2823) );
  DLY4X1 U8437 ( .A(n1133), .Y(n8013) );
  NAND2XL U8438 ( .A(\buff[35][5] ), .B(n9687), .Y(n1133) );
  DLY4X1 U8439 ( .A(n2824), .Y(n8014) );
  OAI221X2 U8440 ( .A0(n1136), .A1(n1108), .B0(n9687), .B1(n9626), .C0(n8015), 
        .Y(n2824) );
  DLY4X1 U8441 ( .A(n1137), .Y(n8015) );
  NAND2XL U8442 ( .A(\buff[35][6] ), .B(n9687), .Y(n1137) );
  DLY4X1 U8443 ( .A(n2825), .Y(n8016) );
  OAI221X2 U8444 ( .A0(n1140), .A1(n1108), .B0(n9687), .B1(n9620), .C0(n8017), 
        .Y(n2825) );
  DLY4X1 U8445 ( .A(n1141), .Y(n8017) );
  NAND2XL U8446 ( .A(\buff[35][7] ), .B(n9687), .Y(n1141) );
  DLY4X1 U8447 ( .A(n2946), .Y(n8018) );
  OAI221XL U8448 ( .A0(n1737), .A1(n1738), .B0(n9686), .B1(n9655), .C0(n8019), 
        .Y(n2946) );
  DLY4X1 U8449 ( .A(n1740), .Y(n8019) );
  NAND2XL U8450 ( .A(\buff[19][0] ), .B(n9686), .Y(n1740) );
  DLY4X1 U8451 ( .A(n2947), .Y(n8020) );
  OAI221X2 U8452 ( .A0(n1746), .A1(n1738), .B0(n9686), .B1(n9648), .C0(n8021), 
        .Y(n2947) );
  DLY4X1 U8453 ( .A(n1747), .Y(n8021) );
  NAND2XL U8454 ( .A(\buff[19][1] ), .B(n9686), .Y(n1747) );
  DLY4X1 U8455 ( .A(n2948), .Y(n8022) );
  OAI221X2 U8456 ( .A0(n1750), .A1(n1738), .B0(n9686), .B1(n9642), .C0(n8023), 
        .Y(n2948) );
  DLY4X1 U8457 ( .A(n1751), .Y(n8023) );
  NAND2XL U8458 ( .A(\buff[19][2] ), .B(n9686), .Y(n1751) );
  DLY4X1 U8459 ( .A(n2949), .Y(n8024) );
  OAI221X2 U8460 ( .A0(n1754), .A1(n1738), .B0(n9686), .B1(n9639), .C0(n8025), 
        .Y(n2949) );
  DLY4X1 U8461 ( .A(n1755), .Y(n8025) );
  NAND2XL U8462 ( .A(\buff[19][3] ), .B(n9686), .Y(n1755) );
  DLY4X1 U8463 ( .A(n2832), .Y(n8026) );
  OAI221X2 U8464 ( .A0(n1175), .A1(n1147), .B0(n9714), .B1(n9626), .C0(n8027), 
        .Y(n2832) );
  DLY4X1 U8465 ( .A(n1176), .Y(n8027) );
  NAND2XL U8466 ( .A(\buff[34][6] ), .B(n9714), .Y(n1176) );
  DLY4X1 U8467 ( .A(n2833), .Y(n8028) );
  OAI221X2 U8468 ( .A0(n1179), .A1(n1147), .B0(n9714), .B1(n9620), .C0(n8029), 
        .Y(n2833) );
  DLY4X1 U8469 ( .A(n1180), .Y(n8029) );
  NAND2XL U8470 ( .A(\buff[34][7] ), .B(n9714), .Y(n1180) );
  DLY4X1 U8471 ( .A(n2954), .Y(n8030) );
  DLY4X1 U8472 ( .A(n1779), .Y(n8031) );
  NAND2XL U8473 ( .A(\buff[18][0] ), .B(n9712), .Y(n1779) );
  OAI221X4 U8474 ( .A0(n1785), .A1(n1777), .B0(n9712), .B1(n9648), .C0(n8032), 
        .Y(n2955) );
  DLY4X1 U8475 ( .A(n8033), .Y(n8032) );
  DLY4X1 U8476 ( .A(n1786), .Y(n8033) );
  NAND2XL U8477 ( .A(\buff[18][1] ), .B(n9712), .Y(n1786) );
  OAI221X4 U8478 ( .A0(n1789), .A1(n1777), .B0(n9712), .B1(n9642), .C0(n8034), 
        .Y(n2956) );
  DLY4X1 U8479 ( .A(n8035), .Y(n8034) );
  DLY4X1 U8480 ( .A(n1790), .Y(n8035) );
  NAND2XL U8481 ( .A(\buff[18][2] ), .B(n9712), .Y(n1790) );
  OAI221X4 U8482 ( .A0(n1793), .A1(n1777), .B0(n9712), .B1(n9639), .C0(n8036), 
        .Y(n2957) );
  DLY4X1 U8483 ( .A(n8037), .Y(n8036) );
  DLY4X1 U8484 ( .A(n1794), .Y(n8037) );
  NAND2XL U8485 ( .A(\buff[18][3] ), .B(n9712), .Y(n1794) );
  OAI221X4 U8486 ( .A0(n1797), .A1(n1777), .B0(n9712), .B1(n9634), .C0(n8038), 
        .Y(n2958) );
  DLY4X1 U8487 ( .A(n8039), .Y(n8038) );
  DLY4X1 U8488 ( .A(n1798), .Y(n8039) );
  NAND2XL U8489 ( .A(\buff[18][4] ), .B(n9712), .Y(n1798) );
  OAI221X4 U8490 ( .A0(n1801), .A1(n1777), .B0(n9712), .B1(n9628), .C0(n8040), 
        .Y(n2959) );
  DLY4X1 U8491 ( .A(n8041), .Y(n8040) );
  DLY4X1 U8492 ( .A(n1802), .Y(n8041) );
  NAND2XL U8493 ( .A(\buff[18][5] ), .B(n9712), .Y(n1802) );
  DLY4X1 U8494 ( .A(n8043), .Y(n8042) );
  DLY4X1 U8495 ( .A(n1532), .Y(n8043) );
  NAND2XL U8496 ( .A(\buff[25][6] ), .B(n9680), .Y(n1532) );
  DLY4X1 U8497 ( .A(n8045), .Y(n8044) );
  DLY4X1 U8498 ( .A(n1536), .Y(n8045) );
  NAND2XL U8499 ( .A(\buff[25][7] ), .B(n9680), .Y(n1536) );
  DLY4X1 U8500 ( .A(n2962), .Y(n8046) );
  DLY4X1 U8501 ( .A(n1820), .Y(n8047) );
  NAND2XL U8502 ( .A(\buff[17][0] ), .B(n9679), .Y(n1820) );
  DLY4X1 U8503 ( .A(n2963), .Y(n8048) );
  DLY4X1 U8504 ( .A(n1827), .Y(n8049) );
  NAND2XL U8505 ( .A(\buff[17][1] ), .B(n9679), .Y(n1827) );
  DLY4X1 U8506 ( .A(n2964), .Y(n8050) );
  DLY4X1 U8507 ( .A(n1831), .Y(n8051) );
  NAND2XL U8508 ( .A(\buff[17][2] ), .B(n9679), .Y(n1831) );
  DLY4X1 U8509 ( .A(n2965), .Y(n8052) );
  DLY4X1 U8510 ( .A(n1835), .Y(n8053) );
  NAND2XL U8511 ( .A(\buff[17][3] ), .B(n9679), .Y(n1835) );
  DLY4X1 U8512 ( .A(n2966), .Y(n8054) );
  DLY4X1 U8513 ( .A(n1839), .Y(n8055) );
  NAND2XL U8514 ( .A(\buff[17][4] ), .B(n9679), .Y(n1839) );
  DLY4X1 U8515 ( .A(n2967), .Y(n8056) );
  DLY4X1 U8516 ( .A(n1843), .Y(n8057) );
  NAND2XL U8517 ( .A(\buff[17][5] ), .B(n9679), .Y(n1843) );
  DLY4X1 U8518 ( .A(n2848), .Y(n8058) );
  OAI221X2 U8519 ( .A0(n1253), .A1(n1225), .B0(n9674), .B1(n9626), .C0(n8059), 
        .Y(n2848) );
  DLY4X1 U8520 ( .A(n1254), .Y(n8059) );
  NAND2XL U8521 ( .A(\buff[32][6] ), .B(n9674), .Y(n1254) );
  DLY4X1 U8522 ( .A(n2849), .Y(n8060) );
  OAI221X2 U8523 ( .A0(n1257), .A1(n1225), .B0(n9674), .B1(n9620), .C0(n8061), 
        .Y(n2849) );
  DLY4X1 U8524 ( .A(n1258), .Y(n8061) );
  NAND2XL U8525 ( .A(\buff[32][7] ), .B(n9674), .Y(n1258) );
  DLY4X1 U8526 ( .A(n2970), .Y(n8062) );
  DLY4X1 U8527 ( .A(n1859), .Y(n8063) );
  NAND2XL U8528 ( .A(\buff[16][0] ), .B(n9672), .Y(n1859) );
  DLY4X1 U8529 ( .A(n2971), .Y(n8064) );
  DLY4X1 U8530 ( .A(n1866), .Y(n8065) );
  NAND2XL U8531 ( .A(\buff[16][1] ), .B(n9672), .Y(n1866) );
  DLY4X1 U8532 ( .A(n2972), .Y(n8066) );
  DLY4X1 U8533 ( .A(n1870), .Y(n8067) );
  NAND2XL U8534 ( .A(\buff[16][2] ), .B(n9672), .Y(n1870) );
  DLY4X1 U8535 ( .A(n2973), .Y(n8068) );
  DLY4X1 U8536 ( .A(n1874), .Y(n8069) );
  NAND2XL U8537 ( .A(\buff[16][3] ), .B(n9672), .Y(n1874) );
  DLY4X1 U8538 ( .A(n2974), .Y(n8070) );
  DLY4X1 U8539 ( .A(n1878), .Y(n8071) );
  NAND2XL U8540 ( .A(\buff[16][4] ), .B(n9672), .Y(n1878) );
  DLY4X1 U8541 ( .A(n2975), .Y(n8072) );
  DLY4X1 U8542 ( .A(n1882), .Y(n8073) );
  NAND2XL U8543 ( .A(\buff[16][5] ), .B(n9672), .Y(n1882) );
  DLY4X1 U8544 ( .A(\buff[31][4] ), .Y(n8074) );
  OAI211XL U8545 ( .A0(n9403), .A1(n9635), .B0(n1284), .C0(n1285), .Y(n2854)
         );
  NAND2XL U8546 ( .A(n8074), .B(n9403), .Y(n1285) );
  DLY4X1 U8547 ( .A(\buff[31][5] ), .Y(n8076) );
  OAI211XL U8548 ( .A0(n9403), .A1(n9628), .B0(n1288), .C0(n1289), .Y(n2855)
         );
  NAND2XL U8549 ( .A(n8076), .B(n9403), .Y(n1289) );
  DLY3X1 U8550 ( .A(n2856), .Y(n8078) );
  OAI211X1 U8551 ( .A0(n9403), .A1(n9624), .B0(n1292), .C0(n8079), .Y(n2856)
         );
  DLY4X1 U8552 ( .A(n1293), .Y(n8079) );
  NAND2XL U8553 ( .A(\buff[31][6] ), .B(n9403), .Y(n1293) );
  DLY4X1 U8554 ( .A(\buff[31][7] ), .Y(n8080) );
  OAI211XL U8555 ( .A0(n9403), .A1(n288), .B0(n1296), .C0(n1297), .Y(n2857) );
  NAND2XL U8556 ( .A(n8080), .B(n9403), .Y(n1297) );
  DLY4X1 U8557 ( .A(n8083), .Y(n8082) );
  OAI211XL U8558 ( .A0(n9383), .A1(n9656), .B0(n1896), .C0(n1897), .Y(n2978)
         );
  NAND2XL U8559 ( .A(\buff[15][0] ), .B(n9383), .Y(n1897) );
  DLY4X1 U8560 ( .A(n8085), .Y(n8084) );
  OAI211XL U8561 ( .A0(n9383), .A1(n9648), .B0(n1904), .C0(n1905), .Y(n2979)
         );
  NAND2XL U8562 ( .A(\buff[15][1] ), .B(n9383), .Y(n1905) );
  DLY4X1 U8563 ( .A(n8087), .Y(n8086) );
  OAI211XL U8564 ( .A0(n9383), .A1(n9642), .B0(n1908), .C0(n1909), .Y(n2980)
         );
  NAND2XL U8565 ( .A(\buff[15][2] ), .B(n9383), .Y(n1909) );
  DLY4X1 U8566 ( .A(n8089), .Y(n8088) );
  OAI211XL U8567 ( .A0(n9383), .A1(n9639), .B0(n1912), .C0(n1913), .Y(n2981)
         );
  NAND2XL U8568 ( .A(\buff[15][3] ), .B(n9383), .Y(n1913) );
  DLY4X1 U8569 ( .A(n8091), .Y(n8090) );
  DLY4X1 U8570 ( .A(n1648), .Y(n8091) );
  NAND2XL U8571 ( .A(\buff[22][6] ), .B(n9705), .Y(n1648) );
  DLY4X1 U8572 ( .A(n8093), .Y(n8092) );
  DLY4X1 U8573 ( .A(n1652), .Y(n8093) );
  NAND2XL U8574 ( .A(\buff[22][7] ), .B(n9705), .Y(n1652) );
  DLY4X1 U8575 ( .A(n8095), .Y(n8094) );
  OAI211XL U8576 ( .A0(n9654), .A1(n9382), .B0(n1935), .C0(n1936), .Y(n2986)
         );
  NAND2XL U8577 ( .A(\buff[14][0] ), .B(n9382), .Y(n1936) );
  DLY4X1 U8578 ( .A(n8097), .Y(n8096) );
  OAI211XL U8579 ( .A0(n9649), .A1(n9382), .B0(n1943), .C0(n1944), .Y(n2987)
         );
  NAND2XL U8580 ( .A(\buff[14][1] ), .B(n9382), .Y(n1944) );
  DLY4X1 U8581 ( .A(n8099), .Y(n8098) );
  OAI211XL U8582 ( .A0(n9643), .A1(n9382), .B0(n1947), .C0(n1948), .Y(n2988)
         );
  NAND2XL U8583 ( .A(\buff[14][2] ), .B(n9382), .Y(n1948) );
  DLY4X1 U8584 ( .A(n8101), .Y(n8100) );
  OAI211XL U8585 ( .A0(n9640), .A1(n9382), .B0(n1951), .C0(n1952), .Y(n2989)
         );
  NAND2XL U8586 ( .A(\buff[14][3] ), .B(n9382), .Y(n1952) );
  DLY4X1 U8587 ( .A(n8103), .Y(n8102) );
  OAI211XL U8588 ( .A0(n9633), .A1(n9382), .B0(n1955), .C0(n1956), .Y(n2990)
         );
  NAND2XL U8589 ( .A(\buff[14][4] ), .B(n9382), .Y(n1956) );
  DLY4X1 U8590 ( .A(n1960), .Y(n8104) );
  DLY4X4 U8591 ( .A(n2991), .Y(n8105) );
  OAI211XL U8592 ( .A0(n9627), .A1(n9382), .B0(n1959), .C0(n8104), .Y(n2991)
         );
  NAND2XL U8593 ( .A(\buff[14][5] ), .B(n9382), .Y(n1960) );
  NAND3X1 U8594 ( .A(n2587), .B(N1657), .C(n2291), .Y(n160) );
  DLY4X1 U8595 ( .A(n8108), .Y(n8107) );
  OAI221X4 U8596 ( .A0(n1688), .A1(n1660), .B0(n9699), .B1(n9625), .C0(n8107), 
        .Y(n2936) );
  DLY4X1 U8597 ( .A(n1689), .Y(n8108) );
  NAND2XL U8598 ( .A(\buff[21][6] ), .B(n9699), .Y(n1689) );
  DLY4X1 U8599 ( .A(n2937), .Y(n8109) );
  OAI221X2 U8600 ( .A0(n1692), .A1(n1660), .B0(n9699), .B1(n9619), .C0(n8110), 
        .Y(n2937) );
  DLY4X1 U8601 ( .A(n1693), .Y(n8110) );
  NAND2XL U8602 ( .A(\buff[21][7] ), .B(n9699), .Y(n1693) );
  DLY4X1 U8603 ( .A(n2994), .Y(n8111) );
  DLY4X1 U8604 ( .A(n1979), .Y(n8112) );
  NAND2XL U8605 ( .A(\buff[13][0] ), .B(n9698), .Y(n1979) );
  OAI221X4 U8606 ( .A0(n1985), .A1(n7224), .B0(n9698), .B1(n9649), .C0(n8113), 
        .Y(n2995) );
  DLY4X1 U8607 ( .A(n8114), .Y(n8113) );
  DLY4X1 U8608 ( .A(n1986), .Y(n8114) );
  NAND2XL U8609 ( .A(\buff[13][1] ), .B(n9698), .Y(n1986) );
  OAI221X4 U8610 ( .A0(n1989), .A1(n7224), .B0(n9698), .B1(n9643), .C0(n8115), 
        .Y(n2996) );
  DLY4X1 U8611 ( .A(n8116), .Y(n8115) );
  DLY4X1 U8612 ( .A(n1990), .Y(n8116) );
  NAND2XL U8613 ( .A(\buff[13][2] ), .B(n9698), .Y(n1990) );
  OAI221X4 U8614 ( .A0(n1993), .A1(n7224), .B0(n9698), .B1(n9640), .C0(n8117), 
        .Y(n2997) );
  DLY4X1 U8615 ( .A(n8118), .Y(n8117) );
  DLY4X1 U8616 ( .A(n1994), .Y(n8118) );
  NAND2XL U8617 ( .A(\buff[13][3] ), .B(n9698), .Y(n1994) );
  OAI221X4 U8618 ( .A0(n1997), .A1(n7224), .B0(n9698), .B1(n9633), .C0(n8119), 
        .Y(n2998) );
  DLY4X1 U8619 ( .A(n8120), .Y(n8119) );
  DLY4X1 U8620 ( .A(n1998), .Y(n8120) );
  NAND2XL U8621 ( .A(\buff[13][4] ), .B(n9698), .Y(n1998) );
  OAI221X4 U8622 ( .A0(n2001), .A1(n7224), .B0(n9698), .B1(n9627), .C0(n8121), 
        .Y(n2999) );
  DLY4X1 U8623 ( .A(n8122), .Y(n8121) );
  DLY4X1 U8624 ( .A(n2002), .Y(n8122) );
  NAND2XL U8625 ( .A(\buff[13][5] ), .B(n9698), .Y(n2002) );
  DLY4X1 U8626 ( .A(n8124), .Y(n8123) );
  DLY4X1 U8627 ( .A(n1728), .Y(n8124) );
  NAND2XL U8628 ( .A(\buff[20][6] ), .B(n9692), .Y(n1728) );
  DLY4X1 U8629 ( .A(n8126), .Y(n8125) );
  DLY4X1 U8630 ( .A(n1732), .Y(n8126) );
  NAND2XL U8631 ( .A(\buff[20][7] ), .B(n9692), .Y(n1732) );
  DLY4X1 U8632 ( .A(n3002), .Y(n8127) );
  DLY4X1 U8633 ( .A(n2018), .Y(n8128) );
  NAND2XL U8634 ( .A(\buff[12][0] ), .B(n9691), .Y(n2018) );
  DLY4X1 U8635 ( .A(n3003), .Y(n8129) );
  DLY4X1 U8636 ( .A(n2025), .Y(n8130) );
  NAND2XL U8637 ( .A(\buff[12][1] ), .B(n9691), .Y(n2025) );
  DLY4X1 U8638 ( .A(n3004), .Y(n8131) );
  DLY4X1 U8639 ( .A(n2029), .Y(n8132) );
  NAND2XL U8640 ( .A(\buff[12][2] ), .B(n9691), .Y(n2029) );
  DLY4X1 U8641 ( .A(n3005), .Y(n8133) );
  DLY4X1 U8642 ( .A(n2033), .Y(n8134) );
  NAND2XL U8643 ( .A(\buff[12][3] ), .B(n9691), .Y(n2033) );
  DLY4X1 U8644 ( .A(n3006), .Y(n8135) );
  DLY4X1 U8645 ( .A(n2037), .Y(n8136) );
  NAND2XL U8646 ( .A(\buff[12][4] ), .B(n9691), .Y(n2037) );
  DLY4X1 U8647 ( .A(n3007), .Y(n8137) );
  DLY4X1 U8648 ( .A(n2041), .Y(n8138) );
  NAND2XL U8649 ( .A(\buff[12][5] ), .B(n9691), .Y(n2041) );
  DLY4X1 U8650 ( .A(n2950), .Y(n8139) );
  OAI221X2 U8651 ( .A0(n1758), .A1(n1738), .B0(n9686), .B1(n9634), .C0(n8140), 
        .Y(n2950) );
  DLY4X1 U8652 ( .A(n1759), .Y(n8140) );
  NAND2XL U8653 ( .A(\buff[19][4] ), .B(n9686), .Y(n1759) );
  DLY4X1 U8654 ( .A(n2951), .Y(n8141) );
  OAI221X2 U8655 ( .A0(n1762), .A1(n1738), .B0(n9686), .B1(n9628), .C0(n8142), 
        .Y(n2951) );
  DLY4X1 U8656 ( .A(n1763), .Y(n8142) );
  NAND2XL U8657 ( .A(\buff[19][5] ), .B(n9686), .Y(n1763) );
  DLY3X4 U8658 ( .A(n2952), .Y(n8143) );
  OAI221X2 U8659 ( .A0(n1766), .A1(n1738), .B0(n9686), .B1(n9624), .C0(n8144), 
        .Y(n2952) );
  DLY4X1 U8660 ( .A(n1767), .Y(n8144) );
  NAND2XL U8661 ( .A(\buff[19][6] ), .B(n9686), .Y(n1767) );
  DLY4X1 U8662 ( .A(n2953), .Y(n8145) );
  OAI221X2 U8663 ( .A0(n1770), .A1(n1738), .B0(n9686), .B1(n9619), .C0(n8146), 
        .Y(n2953) );
  DLY4X1 U8664 ( .A(n1771), .Y(n8146) );
  NAND2XL U8665 ( .A(\buff[19][7] ), .B(n9686), .Y(n1771) );
  DLY4X1 U8666 ( .A(n3010), .Y(n8147) );
  OAI221XL U8667 ( .A0(n2054), .A1(n2055), .B0(n9685), .B1(n9655), .C0(n8148), 
        .Y(n3010) );
  DLY4X1 U8668 ( .A(n2057), .Y(n8148) );
  NAND2XL U8669 ( .A(\buff[11][0] ), .B(n9685), .Y(n2057) );
  DLY4X1 U8670 ( .A(n3011), .Y(n8149) );
  OAI221X2 U8671 ( .A0(n2063), .A1(n2055), .B0(n9685), .B1(n9648), .C0(n8150), 
        .Y(n3011) );
  DLY4X1 U8672 ( .A(n2064), .Y(n8150) );
  NAND2XL U8673 ( .A(\buff[11][1] ), .B(n9685), .Y(n2064) );
  DLY4X1 U8674 ( .A(n3012), .Y(n8151) );
  OAI221X2 U8675 ( .A0(n2067), .A1(n2055), .B0(n9685), .B1(n9642), .C0(n8152), 
        .Y(n3012) );
  DLY4X1 U8676 ( .A(n2068), .Y(n8152) );
  NAND2XL U8677 ( .A(\buff[11][2] ), .B(n9685), .Y(n2068) );
  DLY4X1 U8678 ( .A(n3013), .Y(n8153) );
  OAI221X2 U8679 ( .A0(n2071), .A1(n2055), .B0(n9685), .B1(n9639), .C0(n8154), 
        .Y(n3013) );
  DLY4X1 U8680 ( .A(n2072), .Y(n8154) );
  NAND2XL U8681 ( .A(\buff[11][3] ), .B(n9685), .Y(n2072) );
  OAI221X4 U8682 ( .A0(n1805), .A1(n1777), .B0(n9712), .B1(n9624), .C0(n8155), 
        .Y(n2960) );
  DLY4X1 U8683 ( .A(n8156), .Y(n8155) );
  DLY4X1 U8684 ( .A(n1806), .Y(n8156) );
  NAND2XL U8685 ( .A(\buff[18][6] ), .B(n9712), .Y(n1806) );
  OAI221X4 U8686 ( .A0(n1809), .A1(n1777), .B0(n9712), .B1(n9619), .C0(n8157), 
        .Y(n2961) );
  DLY4X1 U8687 ( .A(n8158), .Y(n8157) );
  DLY4X1 U8688 ( .A(n1810), .Y(n8158) );
  NAND2XL U8689 ( .A(\buff[18][7] ), .B(n9712), .Y(n1810) );
  DLY4X1 U8690 ( .A(n3018), .Y(n8159) );
  DLY4X1 U8691 ( .A(n2096), .Y(n8160) );
  NAND2XL U8692 ( .A(\buff[10][0] ), .B(n9711), .Y(n2096) );
  OAI221X4 U8693 ( .A0(n2102), .A1(n2094), .B0(n9711), .B1(n9649), .C0(n8161), 
        .Y(n3019) );
  DLY4X1 U8694 ( .A(n8162), .Y(n8161) );
  DLY4X1 U8695 ( .A(n2103), .Y(n8162) );
  NAND2XL U8696 ( .A(\buff[10][1] ), .B(n9711), .Y(n2103) );
  OAI221X4 U8697 ( .A0(n2106), .A1(n2094), .B0(n9711), .B1(n9643), .C0(n8163), 
        .Y(n3020) );
  DLY4X1 U8698 ( .A(n8164), .Y(n8163) );
  DLY4X1 U8699 ( .A(n2107), .Y(n8164) );
  NAND2XL U8700 ( .A(\buff[10][2] ), .B(n9711), .Y(n2107) );
  OAI221X4 U8701 ( .A0(n2110), .A1(n2094), .B0(n9711), .B1(n9640), .C0(n8165), 
        .Y(n3021) );
  DLY4X1 U8702 ( .A(n8166), .Y(n8165) );
  DLY4X1 U8703 ( .A(n2111), .Y(n8166) );
  NAND2XL U8704 ( .A(\buff[10][3] ), .B(n9711), .Y(n2111) );
  OAI221X4 U8705 ( .A0(n2114), .A1(n2094), .B0(n9711), .B1(n9633), .C0(n8167), 
        .Y(n3022) );
  DLY4X1 U8706 ( .A(n8168), .Y(n8167) );
  DLY4X1 U8707 ( .A(n2115), .Y(n8168) );
  NAND2XL U8708 ( .A(\buff[10][4] ), .B(n9711), .Y(n2115) );
  OAI221X4 U8709 ( .A0(n2118), .A1(n2094), .B0(n9711), .B1(n9627), .C0(n8169), 
        .Y(n3023) );
  DLY4X1 U8710 ( .A(n8170), .Y(n8169) );
  DLY4X1 U8711 ( .A(n2119), .Y(n8170) );
  NAND2XL U8712 ( .A(\buff[10][5] ), .B(n9711), .Y(n2119) );
  DLY4X1 U8713 ( .A(n8172), .Y(n8171) );
  DLY4X1 U8714 ( .A(n1847), .Y(n8172) );
  NAND2XL U8715 ( .A(\buff[17][6] ), .B(n9679), .Y(n1847) );
  DLY4X1 U8716 ( .A(n8174), .Y(n8173) );
  DLY4X1 U8717 ( .A(n1851), .Y(n8174) );
  NAND2XL U8718 ( .A(\buff[17][7] ), .B(n9679), .Y(n1851) );
  DLY4X1 U8719 ( .A(n3026), .Y(n8175) );
  DLY4X1 U8720 ( .A(n2139), .Y(n8176) );
  NAND2XL U8721 ( .A(\buff[9][0] ), .B(n9678), .Y(n2139) );
  DLY4X1 U8722 ( .A(n3027), .Y(n8177) );
  DLY4X1 U8723 ( .A(n2146), .Y(n8178) );
  NAND2XL U8724 ( .A(\buff[9][1] ), .B(n9678), .Y(n2146) );
  DLY4X1 U8725 ( .A(n3028), .Y(n8179) );
  DLY4X1 U8726 ( .A(n2150), .Y(n8180) );
  NAND2XL U8727 ( .A(\buff[9][2] ), .B(n9678), .Y(n2150) );
  DLY4X1 U8728 ( .A(n3029), .Y(n8181) );
  DLY4X1 U8729 ( .A(n2154), .Y(n8182) );
  NAND2XL U8730 ( .A(\buff[9][3] ), .B(n9678), .Y(n2154) );
  DLY4X1 U8731 ( .A(n3030), .Y(n8183) );
  DLY4X1 U8732 ( .A(n2158), .Y(n8184) );
  NAND2XL U8733 ( .A(\buff[9][4] ), .B(n9678), .Y(n2158) );
  DLY4X1 U8734 ( .A(n3031), .Y(n8185) );
  DLY4X1 U8735 ( .A(n2162), .Y(n8186) );
  NAND2XL U8736 ( .A(\buff[9][5] ), .B(n9678), .Y(n2162) );
  BUFX2 U8737 ( .A(n1654), .Y(n8187) );
  DLY4X1 U8738 ( .A(\buff[16][6] ), .Y(n8188) );
  OAI221X4 U8739 ( .A0(n1885), .A1(n1857), .B0(n9672), .B1(n9624), .C0(n8189), 
        .Y(n2976) );
  DLY4X1 U8740 ( .A(n1886), .Y(n8189) );
  NAND2XL U8741 ( .A(n8188), .B(n9672), .Y(n1886) );
  DLY4X1 U8742 ( .A(n2977), .Y(n8190) );
  OAI221X2 U8743 ( .A0(n1889), .A1(n1857), .B0(n9672), .B1(n9619), .C0(n8191), 
        .Y(n2977) );
  DLY4X1 U8744 ( .A(n1890), .Y(n8191) );
  NAND2XL U8745 ( .A(\buff[16][7] ), .B(n9672), .Y(n1890) );
  DLY4X1 U8746 ( .A(n3034), .Y(n8192) );
  DLY4X1 U8747 ( .A(n2178), .Y(n8193) );
  NAND2XL U8748 ( .A(\buff[8][0] ), .B(n9671), .Y(n2178) );
  DLY4X1 U8749 ( .A(n3035), .Y(n8194) );
  DLY4X1 U8750 ( .A(n2185), .Y(n8195) );
  NAND2XL U8751 ( .A(\buff[8][1] ), .B(n9671), .Y(n2185) );
  DLY4X1 U8752 ( .A(n3036), .Y(n8196) );
  DLY4X1 U8753 ( .A(n2189), .Y(n8197) );
  NAND2XL U8754 ( .A(\buff[8][2] ), .B(n9671), .Y(n2189) );
  DLY4X1 U8755 ( .A(n3037), .Y(n8198) );
  DLY4X1 U8756 ( .A(n2193), .Y(n8199) );
  NAND2XL U8757 ( .A(\buff[8][3] ), .B(n9671), .Y(n2193) );
  DLY4X1 U8758 ( .A(n3038), .Y(n8200) );
  DLY4X1 U8759 ( .A(n2197), .Y(n8201) );
  NAND2XL U8760 ( .A(\buff[8][4] ), .B(n9671), .Y(n2197) );
  DLY4X1 U8761 ( .A(n3039), .Y(n8202) );
  DLY4X1 U8762 ( .A(n2201), .Y(n8203) );
  NAND2XL U8763 ( .A(\buff[8][5] ), .B(n9671), .Y(n2201) );
  DLY4X1 U8764 ( .A(\buff[15][4] ), .Y(n8204) );
  OAI211XL U8765 ( .A0(n9383), .A1(n9635), .B0(n1916), .C0(n1917), .Y(n2982)
         );
  NAND2XL U8766 ( .A(n8204), .B(n9383), .Y(n1917) );
  DLY4X1 U8767 ( .A(\buff[15][5] ), .Y(n8206) );
  OAI211XL U8768 ( .A0(n9383), .A1(n9629), .B0(n1920), .C0(n1921), .Y(n2983)
         );
  NAND2XL U8769 ( .A(n8206), .B(n9383), .Y(n1921) );
  DLY4X1 U8770 ( .A(\buff[15][6] ), .Y(n8208) );
  OAI211XL U8771 ( .A0(n9383), .A1(n9625), .B0(n1924), .C0(n1925), .Y(n2984)
         );
  NAND2XL U8772 ( .A(n8208), .B(n9383), .Y(n1925) );
  DLY4X1 U8773 ( .A(\buff[15][7] ), .Y(n8210) );
  OAI211XL U8774 ( .A0(n9383), .A1(n288), .B0(n1928), .C0(n1929), .Y(n2985) );
  NAND2XL U8775 ( .A(n8210), .B(n9383), .Y(n1929) );
  DLY4X1 U8776 ( .A(n8213), .Y(n8212) );
  OAI211XL U8777 ( .A0(n9375), .A1(n9655), .B0(n2215), .C0(n2216), .Y(n3042)
         );
  NAND2XL U8778 ( .A(\buff[7][0] ), .B(n9375), .Y(n2216) );
  DLY4X1 U8779 ( .A(n8215), .Y(n8214) );
  OAI211XL U8780 ( .A0(n9375), .A1(n9648), .B0(n2223), .C0(n2224), .Y(n3043)
         );
  NAND2XL U8781 ( .A(\buff[7][1] ), .B(n9375), .Y(n2224) );
  DLY4X1 U8782 ( .A(n8217), .Y(n8216) );
  OAI211XL U8783 ( .A0(n9375), .A1(n9642), .B0(n2227), .C0(n2228), .Y(n3044)
         );
  NAND2XL U8784 ( .A(\buff[7][2] ), .B(n9375), .Y(n2228) );
  DLY4X1 U8785 ( .A(n8219), .Y(n8218) );
  OAI211XL U8786 ( .A0(n9375), .A1(n9639), .B0(n2231), .C0(n2232), .Y(n3045)
         );
  NAND2XL U8787 ( .A(\buff[7][3] ), .B(n9375), .Y(n2232) );
  DLY4X1 U8788 ( .A(n8221), .Y(n8220) );
  OAI211X4 U8789 ( .A0(n9625), .A1(n9382), .B0(n1963), .C0(n8220), .Y(n2992)
         );
  DLY4X1 U8790 ( .A(n1964), .Y(n8221) );
  NAND2XL U8791 ( .A(\buff[14][6] ), .B(n9382), .Y(n1964) );
  DLY4X1 U8792 ( .A(n1968), .Y(n8222) );
  DLY4X4 U8793 ( .A(n2993), .Y(n8223) );
  OAI211XL U8794 ( .A0(n9618), .A1(n9382), .B0(n1967), .C0(n8222), .Y(n2993)
         );
  NAND2XL U8795 ( .A(\buff[14][7] ), .B(n9382), .Y(n1968) );
  OAI221X4 U8796 ( .A0(n2254), .A1(n2255), .B0(n9704), .B1(n9654), .C0(n8224), 
        .Y(n3050) );
  DLY4X1 U8797 ( .A(n8225), .Y(n8224) );
  DLY4X1 U8798 ( .A(n2257), .Y(n8225) );
  NAND2XL U8799 ( .A(\buff[6][0] ), .B(n9704), .Y(n2257) );
  OAI221X4 U8800 ( .A0(n2262), .A1(n2255), .B0(n9704), .B1(n9649), .C0(n8226), 
        .Y(n3051) );
  DLY4X1 U8801 ( .A(n8227), .Y(n8226) );
  DLY4X1 U8802 ( .A(n2263), .Y(n8227) );
  NAND2XL U8803 ( .A(\buff[6][1] ), .B(n9704), .Y(n2263) );
  OAI221X4 U8804 ( .A0(n2266), .A1(n2255), .B0(n9704), .B1(n9643), .C0(n8228), 
        .Y(n3052) );
  DLY4X1 U8805 ( .A(n8229), .Y(n8228) );
  DLY4X1 U8806 ( .A(n2267), .Y(n8229) );
  NAND2XL U8807 ( .A(\buff[6][2] ), .B(n9704), .Y(n2267) );
  OAI221X4 U8808 ( .A0(n2270), .A1(n2255), .B0(n9704), .B1(n9640), .C0(n8230), 
        .Y(n3053) );
  DLY4X1 U8809 ( .A(n8231), .Y(n8230) );
  DLY4X1 U8810 ( .A(n2271), .Y(n8231) );
  NAND2XL U8811 ( .A(\buff[6][3] ), .B(n9704), .Y(n2271) );
  OAI221X4 U8812 ( .A0(n2274), .A1(n2255), .B0(n9704), .B1(n9633), .C0(n8232), 
        .Y(n3054) );
  DLY4X1 U8813 ( .A(n8233), .Y(n8232) );
  DLY4X1 U8814 ( .A(n2275), .Y(n8233) );
  NAND2XL U8815 ( .A(\buff[6][4] ), .B(n9704), .Y(n2275) );
  OAI221X4 U8816 ( .A0(n2278), .A1(n2255), .B0(n9704), .B1(n9627), .C0(n8234), 
        .Y(n3055) );
  DLY4X1 U8817 ( .A(n8235), .Y(n8234) );
  DLY4X1 U8818 ( .A(n2279), .Y(n8235) );
  NAND2XL U8819 ( .A(\buff[6][5] ), .B(n9704), .Y(n2279) );
  DLY4X1 U8820 ( .A(n3000), .Y(n8236) );
  OAI221X2 U8821 ( .A0(n2005), .A1(n1977), .B0(n9698), .B1(n9625), .C0(n8237), 
        .Y(n3000) );
  DLY4X1 U8822 ( .A(n2006), .Y(n8237) );
  NAND2XL U8823 ( .A(\buff[13][6] ), .B(n9698), .Y(n2006) );
  DLY4X1 U8824 ( .A(n3001), .Y(n8238) );
  OAI221X2 U8825 ( .A0(n2009), .A1(n1977), .B0(n9698), .B1(n9618), .C0(n8239), 
        .Y(n3001) );
  DLY4X1 U8826 ( .A(n2010), .Y(n8239) );
  NAND2XL U8827 ( .A(\buff[13][7] ), .B(n9698), .Y(n2010) );
  DLY4X1 U8828 ( .A(n3058), .Y(n8240) );
  DLY4X1 U8829 ( .A(n2298), .Y(n8241) );
  NAND2XL U8830 ( .A(\buff[5][0] ), .B(n9697), .Y(n2298) );
  DLY4X1 U8831 ( .A(n3059), .Y(n8242) );
  DLY4X1 U8832 ( .A(n2306), .Y(n8243) );
  NAND2XL U8833 ( .A(\buff[5][1] ), .B(n9697), .Y(n2306) );
  DLY4X1 U8834 ( .A(n3060), .Y(n8244) );
  DLY4X1 U8835 ( .A(n2310), .Y(n8245) );
  NAND2XL U8836 ( .A(\buff[5][2] ), .B(n9697), .Y(n2310) );
  DLY4X1 U8837 ( .A(n3061), .Y(n8246) );
  DLY4X1 U8838 ( .A(n2314), .Y(n8247) );
  NAND2XL U8839 ( .A(\buff[5][3] ), .B(n9697), .Y(n2314) );
  NAND2XL U8840 ( .A(n9661), .B(n2331), .Y(n2296) );
  BUFX2 U8841 ( .A(n2296), .Y(n8248) );
  OAI221X4 U8842 ( .A0(n2317), .A1(n8248), .B0(n9697), .B1(n9633), .C0(n8249), 
        .Y(n3062) );
  DLY4X1 U8843 ( .A(n8250), .Y(n8249) );
  DLY4X1 U8844 ( .A(n2318), .Y(n8250) );
  NAND2XL U8845 ( .A(\buff[5][4] ), .B(n9697), .Y(n2318) );
  DLY4X1 U8846 ( .A(n3063), .Y(n8251) );
  OAI221X2 U8847 ( .A0(n2321), .A1(n2296), .B0(n9697), .B1(n9627), .C0(n8252), 
        .Y(n3063) );
  DLY4X1 U8848 ( .A(n2322), .Y(n8252) );
  NAND2XL U8849 ( .A(\buff[5][5] ), .B(n9697), .Y(n2322) );
  DLY4X1 U8850 ( .A(n8254), .Y(n8253) );
  DLY4X1 U8851 ( .A(n2045), .Y(n8254) );
  NAND2XL U8852 ( .A(\buff[12][6] ), .B(n9691), .Y(n2045) );
  DLY4X1 U8853 ( .A(n8256), .Y(n8255) );
  DLY4X1 U8854 ( .A(n2049), .Y(n8256) );
  NAND2XL U8855 ( .A(\buff[12][7] ), .B(n9691), .Y(n2049) );
  DLY4X1 U8856 ( .A(n3066), .Y(n8257) );
  DLY4X1 U8857 ( .A(n2338), .Y(n8258) );
  NAND2XL U8858 ( .A(\buff[4][0] ), .B(n9690), .Y(n2338) );
  DLY4X1 U8859 ( .A(n3067), .Y(n8259) );
  DLY4X1 U8860 ( .A(n2346), .Y(n8260) );
  NAND2XL U8861 ( .A(\buff[4][1] ), .B(n9690), .Y(n2346) );
  DLY4X1 U8862 ( .A(n3068), .Y(n8261) );
  DLY4X1 U8863 ( .A(n2350), .Y(n8262) );
  NAND2XL U8864 ( .A(\buff[4][2] ), .B(n9690), .Y(n2350) );
  BUFX2 U8865 ( .A(n173), .Y(n8263) );
  OAI221X4 U8866 ( .A0(n2353), .A1(n2336), .B0(n9690), .B1(n9640), .C0(n8264), 
        .Y(n3069) );
  DLY4X1 U8867 ( .A(n8265), .Y(n8264) );
  DLY4X1 U8868 ( .A(n2354), .Y(n8265) );
  NAND2XL U8869 ( .A(\buff[4][3] ), .B(n9690), .Y(n2354) );
  DLY4X1 U8870 ( .A(n3070), .Y(n8266) );
  OAI221X2 U8871 ( .A0(n2357), .A1(n2336), .B0(n9690), .B1(n9633), .C0(n8267), 
        .Y(n3070) );
  DLY4X1 U8872 ( .A(n2358), .Y(n8267) );
  NAND2XL U8873 ( .A(\buff[4][4] ), .B(n9690), .Y(n2358) );
  DLY4X1 U8874 ( .A(n3071), .Y(n8268) );
  OAI221X2 U8875 ( .A0(n2361), .A1(n2336), .B0(n9690), .B1(n9627), .C0(n8269), 
        .Y(n3071) );
  DLY4X1 U8876 ( .A(n2362), .Y(n8269) );
  NAND2XL U8877 ( .A(\buff[4][5] ), .B(n9690), .Y(n2362) );
  DLY4X1 U8878 ( .A(n3014), .Y(n8270) );
  OAI221X2 U8879 ( .A0(n2075), .A1(n2055), .B0(n9685), .B1(n9634), .C0(n8271), 
        .Y(n3014) );
  DLY4X1 U8880 ( .A(n2076), .Y(n8271) );
  NAND2XL U8881 ( .A(\buff[11][4] ), .B(n9685), .Y(n2076) );
  DLY4X1 U8882 ( .A(n3015), .Y(n8272) );
  OAI221X2 U8883 ( .A0(n2079), .A1(n2055), .B0(n9685), .B1(n9628), .C0(n8273), 
        .Y(n3015) );
  DLY4X1 U8884 ( .A(n2080), .Y(n8273) );
  NAND2XL U8885 ( .A(\buff[11][5] ), .B(n9685), .Y(n2080) );
  DLY4X1 U8886 ( .A(n3016), .Y(n8274) );
  OAI221X2 U8887 ( .A0(n2083), .A1(n2055), .B0(n9685), .B1(n9626), .C0(n8275), 
        .Y(n3016) );
  DLY4X1 U8888 ( .A(n2084), .Y(n8275) );
  NAND2XL U8889 ( .A(\buff[11][6] ), .B(n9685), .Y(n2084) );
  DLY4X1 U8890 ( .A(n3017), .Y(n8276) );
  OAI221X2 U8891 ( .A0(n2087), .A1(n2055), .B0(n9685), .B1(n9619), .C0(n8277), 
        .Y(n3017) );
  DLY4X1 U8892 ( .A(n2088), .Y(n8277) );
  NAND2XL U8893 ( .A(\buff[11][7] ), .B(n9685), .Y(n2088) );
  DLY4X1 U8894 ( .A(n3074), .Y(n8278) );
  OAI221X2 U8895 ( .A0(n2375), .A1(n2376), .B0(n9684), .B1(n9655), .C0(n8279), 
        .Y(n3074) );
  DLY4X1 U8896 ( .A(n2378), .Y(n8279) );
  NAND2XL U8897 ( .A(\buff[3][0] ), .B(n9684), .Y(n2378) );
  DLY4X1 U8898 ( .A(n3075), .Y(n8280) );
  OAI221X2 U8899 ( .A0(n2385), .A1(n2376), .B0(n9684), .B1(n9648), .C0(n8281), 
        .Y(n3075) );
  DLY4X1 U8900 ( .A(n2386), .Y(n8281) );
  NAND2XL U8901 ( .A(\buff[3][1] ), .B(n9684), .Y(n2386) );
  DLY4X1 U8902 ( .A(n3076), .Y(n8282) );
  OAI221X2 U8903 ( .A0(n2389), .A1(n2376), .B0(n9684), .B1(n9642), .C0(n8283), 
        .Y(n3076) );
  DLY4X1 U8904 ( .A(n2390), .Y(n8283) );
  NAND2XL U8905 ( .A(\buff[3][2] ), .B(n9684), .Y(n2390) );
  DLY4X1 U8906 ( .A(n3077), .Y(n8284) );
  OAI221X2 U8907 ( .A0(n2393), .A1(n2376), .B0(n9684), .B1(n9639), .C0(n8285), 
        .Y(n3077) );
  DLY4X1 U8908 ( .A(n2394), .Y(n8285) );
  NAND2XL U8909 ( .A(\buff[3][3] ), .B(n9684), .Y(n2394) );
  OAI221X4 U8910 ( .A0(n2122), .A1(n2094), .B0(n9711), .B1(n9625), .C0(n8286), 
        .Y(n3024) );
  DLY4X1 U8911 ( .A(n8287), .Y(n8286) );
  DLY4X1 U8912 ( .A(n2123), .Y(n8287) );
  NAND2XL U8913 ( .A(\buff[10][6] ), .B(n9711), .Y(n2123) );
  OAI221X4 U8914 ( .A0(n2126), .A1(n2094), .B0(n9711), .B1(n9618), .C0(n8288), 
        .Y(n3025) );
  DLY4X1 U8915 ( .A(n8289), .Y(n8288) );
  DLY4X1 U8916 ( .A(n2127), .Y(n8289) );
  NAND2XL U8917 ( .A(\buff[10][7] ), .B(n9711), .Y(n2127) );
  DLY4X1 U8918 ( .A(\buff[2][0] ), .Y(n8290) );
  OAI211XL U8919 ( .A0(n9654), .A1(n9360), .B0(n2416), .C0(n2417), .Y(n3082)
         );
  NAND2XL U8920 ( .A(n8290), .B(n9360), .Y(n2417) );
  DLY4X1 U8921 ( .A(\buff[2][1] ), .Y(n8292) );
  OAI211XL U8922 ( .A0(n9649), .A1(n9360), .B0(n2424), .C0(n2425), .Y(n3083)
         );
  NAND2XL U8923 ( .A(n8292), .B(n9360), .Y(n2425) );
  DLY4X1 U8924 ( .A(\buff[2][2] ), .Y(n8294) );
  OAI211XL U8925 ( .A0(n9643), .A1(n9360), .B0(n2428), .C0(n2429), .Y(n3084)
         );
  NAND2XL U8926 ( .A(n8294), .B(n9360), .Y(n2429) );
  DLY4X1 U8927 ( .A(\buff[2][3] ), .Y(n8296) );
  OAI211XL U8928 ( .A0(n9640), .A1(n9360), .B0(n2432), .C0(n2433), .Y(n3085)
         );
  NAND2XL U8929 ( .A(n8296), .B(n9360), .Y(n2433) );
  DLY4X1 U8930 ( .A(\buff[2][4] ), .Y(n8298) );
  OAI211XL U8931 ( .A0(n9633), .A1(n9360), .B0(n2436), .C0(n2437), .Y(n3086)
         );
  NAND2XL U8932 ( .A(n8298), .B(n9360), .Y(n2437) );
  DLY4X1 U8933 ( .A(\buff[2][5] ), .Y(n8300) );
  OAI211XL U8934 ( .A0(n9627), .A1(n9360), .B0(n2440), .C0(n2441), .Y(n3087)
         );
  NAND2XL U8935 ( .A(n8300), .B(n9360), .Y(n2441) );
  DLY4X1 U8936 ( .A(n8303), .Y(n8302) );
  DLY4X1 U8937 ( .A(n2166), .Y(n8303) );
  NAND2XL U8938 ( .A(\buff[9][6] ), .B(n9678), .Y(n2166) );
  DLY4X1 U8939 ( .A(n8305), .Y(n8304) );
  DLY4X1 U8940 ( .A(n2170), .Y(n8305) );
  NAND2XL U8941 ( .A(\buff[9][7] ), .B(n9678), .Y(n2170) );
  DLY4X1 U8942 ( .A(n3090), .Y(n8306) );
  DLY4X1 U8943 ( .A(n2458), .Y(n8307) );
  NAND2XL U8944 ( .A(\buff[1][0] ), .B(n9677), .Y(n2458) );
  DLY4X1 U8945 ( .A(n3091), .Y(n8308) );
  DLY4X1 U8946 ( .A(n2465), .Y(n8309) );
  NAND2XL U8947 ( .A(\buff[1][1] ), .B(n9677), .Y(n2465) );
  DLY4X1 U8948 ( .A(n3092), .Y(n8310) );
  DLY4X1 U8949 ( .A(n2469), .Y(n8311) );
  NAND2XL U8950 ( .A(\buff[1][2] ), .B(n9677), .Y(n2469) );
  BUFX2 U8951 ( .A(n212), .Y(n8312) );
  OAI221X4 U8952 ( .A0(n2472), .A1(n2456), .B0(n9677), .B1(n9640), .C0(n8313), 
        .Y(n3093) );
  DLY4X1 U8953 ( .A(n8314), .Y(n8313) );
  DLY4X1 U8954 ( .A(n2473), .Y(n8314) );
  NAND2XL U8955 ( .A(\buff[1][3] ), .B(n9677), .Y(n2473) );
  DLY4X1 U8956 ( .A(n3094), .Y(n8315) );
  OAI221X2 U8957 ( .A0(n2476), .A1(n2456), .B0(n9677), .B1(n9633), .C0(n8316), 
        .Y(n3094) );
  DLY4X1 U8958 ( .A(n2477), .Y(n8316) );
  NAND2XL U8959 ( .A(\buff[1][4] ), .B(n9677), .Y(n2477) );
  DLY4X1 U8960 ( .A(n3095), .Y(n8317) );
  OAI221X2 U8961 ( .A0(n2480), .A1(n2456), .B0(n9677), .B1(n9627), .C0(n8318), 
        .Y(n3095) );
  DLY4X1 U8962 ( .A(n2481), .Y(n8318) );
  NAND2XL U8963 ( .A(\buff[1][5] ), .B(n9677), .Y(n2481) );
  CLKBUFX2 U8964 ( .A(n2582), .Y(n8385) );
  DLY4X1 U8965 ( .A(n8320), .Y(n8319) );
  DLY4X1 U8966 ( .A(n2205), .Y(n8320) );
  NAND2XL U8967 ( .A(\buff[8][6] ), .B(n9671), .Y(n2205) );
  DLY4X1 U8968 ( .A(n3041), .Y(n8321) );
  OAI221X2 U8969 ( .A0(n2208), .A1(n2176), .B0(n9671), .B1(n9618), .C0(n8322), 
        .Y(n3041) );
  DLY4X1 U8970 ( .A(n2209), .Y(n8322) );
  NAND2XL U8971 ( .A(\buff[8][7] ), .B(n9671), .Y(n2209) );
  DLY4X1 U8972 ( .A(n3098), .Y(n8323) );
  DLY4X1 U8973 ( .A(n2497), .Y(n8324) );
  NAND2XL U8974 ( .A(\buff[0][0] ), .B(n9670), .Y(n2497) );
  DLY4X1 U8975 ( .A(n3099), .Y(n8325) );
  DLY4X1 U8976 ( .A(n2506), .Y(n8326) );
  NAND2XL U8977 ( .A(\buff[0][1] ), .B(n9670), .Y(n2506) );
  DLY4X1 U8978 ( .A(n3100), .Y(n8327) );
  DLY4X1 U8979 ( .A(n2510), .Y(n8328) );
  NAND2XL U8980 ( .A(\buff[0][2] ), .B(n9670), .Y(n2510) );
  BUFX2 U8981 ( .A(n227), .Y(n8329) );
  OAI221X4 U8982 ( .A0(n2513), .A1(n2495), .B0(n9670), .B1(n9639), .C0(n8330), 
        .Y(n3101) );
  DLY4X1 U8983 ( .A(n8331), .Y(n8330) );
  DLY4X1 U8984 ( .A(n2514), .Y(n8331) );
  NAND2XL U8985 ( .A(\buff[0][3] ), .B(n9670), .Y(n2514) );
  DLY4X1 U8986 ( .A(n3102), .Y(n8332) );
  OAI221X2 U8987 ( .A0(n2517), .A1(n2495), .B0(n9670), .B1(n9634), .C0(n8333), 
        .Y(n3102) );
  DLY4X1 U8988 ( .A(n2518), .Y(n8333) );
  NAND2XL U8989 ( .A(\buff[0][4] ), .B(n9670), .Y(n2518) );
  DLY4X1 U8990 ( .A(n3103), .Y(n8334) );
  OAI221X2 U8991 ( .A0(n2521), .A1(n2495), .B0(n9670), .B1(n9628), .C0(n8335), 
        .Y(n3103) );
  DLY4X1 U8992 ( .A(n2522), .Y(n8335) );
  NAND2XL U8993 ( .A(\buff[0][5] ), .B(n9670), .Y(n2522) );
  BUFX2 U8994 ( .A(n2601), .Y(n8336) );
  DLY4X4 U8995 ( .A(n8338), .Y(n8337) );
  OAI2BB1XL U8996 ( .A0N(n8337), .A1N(n9458), .B0(n121), .Y(n2601) );
  DLY4X1 U8997 ( .A(n3112), .Y(n8340) );
  BUFX2 U8998 ( .A(n8340), .Y(n8339) );
  OAI21XL U8999 ( .A0(n8372), .A1(n2559), .B0(n2560), .Y(n3112) );
  DLY3X1 U9000 ( .A(n3048), .Y(n8341) );
  OAI211XL U9001 ( .A0(n9375), .A1(n9625), .B0(n2243), .C0(n8342), .Y(n3048)
         );
  DLY4X1 U9002 ( .A(n2244), .Y(n8342) );
  NAND2XL U9003 ( .A(\buff[7][6] ), .B(n9375), .Y(n2244) );
  DLY4X1 U9004 ( .A(n8344), .Y(n8343) );
  DLY4X1 U9005 ( .A(n8346), .Y(n8345) );
  DLY4X1 U9006 ( .A(n8348), .Y(n8347) );
  DLY2X1 U9007 ( .A(next[0]), .Y(n8348) );
  OAI21X4 U9008 ( .A0(n92), .A1(n9665), .B0(n9745), .Y(next[0]) );
  DLY4X1 U9009 ( .A(n8350), .Y(n8349) );
  DLY4X1 U9010 ( .A(n2572), .Y(n8350) );
  NAND2XL U9011 ( .A(n8349), .B(n9745), .Y(n2573) );
  DLY4X1 U9012 ( .A(n2248), .Y(n8352) );
  DLY4X4 U9013 ( .A(n3049), .Y(n8353) );
  OAI211XL U9014 ( .A0(n9375), .A1(n288), .B0(n2247), .C0(n8352), .Y(n3049) );
  NAND2XL U9015 ( .A(\buff[7][7] ), .B(n9375), .Y(n2248) );
  DLY3X1 U9016 ( .A(n2920), .Y(n8354) );
  OAI211XL U9017 ( .A0(n9393), .A1(n9625), .B0(n1609), .C0(n8355), .Y(n2920)
         );
  DLY4X1 U9018 ( .A(n1610), .Y(n8355) );
  NAND2XL U9019 ( .A(\buff[23][6] ), .B(n9393), .Y(n1610) );
  DLY4X1 U9020 ( .A(n8358), .Y(n8357) );
  DLY4X1 U9021 ( .A(\buff[61][6] ), .Y(n8358) );
  BUFX2 U9022 ( .A(n8357), .Y(n8356) );
  DLY4X4 U9023 ( .A(n148), .Y(n9456) );
  DLY4X1 U9024 ( .A(n8360), .Y(n8359) );
  OAI32XL U9025 ( .A0(n2549), .A1(n2550), .A2(n9508), .B0(n2576), .B1(n2551), 
        .Y(n3109) );
  BUFX2 U9026 ( .A(n2600), .Y(n8361) );
  DLY4X4 U9027 ( .A(n8363), .Y(n8362) );
  OAI2BB1XL U9028 ( .A0N(n8362), .A1N(n9458), .B0(n118), .Y(n2600) );
  BUFX2 U9029 ( .A(n8365), .Y(n8364) );
  DLY4X1 U9030 ( .A(n3111), .Y(n8365) );
  CLKBUFX2 U9031 ( .A(n9815), .Y(n9509) );
  INVXL U9032 ( .A(n2575), .Y(n9815) );
  NAND2XL U9033 ( .A(n2571), .B(n9743), .Y(n94) );
  BUFX2 U9034 ( .A(n8367), .Y(n8366) );
  DLY4X4 U9035 ( .A(n8368), .Y(n8367) );
  DLY4X4 U9036 ( .A(n3106), .Y(n8368) );
  OAI32X2 U9037 ( .A0(n2538), .A1(n2539), .A2(n9513), .B0(n9512), .B1(n2540), 
        .Y(n3106) );
  DLY4X1 U9038 ( .A(n3107), .Y(n8369) );
  DLY4X1 U9039 ( .A(n3110), .Y(n8371) );
  DLY4X1 U9040 ( .A(n2588), .Y(n8372) );
  DLY4X4 U9041 ( .A(n8375), .Y(n8374) );
  DLY4X4 U9042 ( .A(n3115), .Y(n8375) );
  DLY4X1 U9043 ( .A(n3117), .Y(n8378) );
  BUFX2 U9044 ( .A(n8377), .Y(n8376) );
  DLY4X1 U9045 ( .A(n8378), .Y(n8377) );
  OAI2BB2X1 U9046 ( .B0(n2586), .B1(n2565), .A0N(N1744), .A1N(n2566), .Y(n3117) );
  DLY4X1 U9047 ( .A(n8381), .Y(n8380) );
  BUFX2 U9048 ( .A(n8380), .Y(n8379) );
  DLY4X1 U9049 ( .A(n3118), .Y(n8381) );
  OAI2BB2X1 U9050 ( .B0(n2587), .B1(n2565), .A0N(N1743), .A1N(n2566), .Y(n3118) );
  BUFX2 U9051 ( .A(n8384), .Y(n8382) );
  DLY4X1 U9052 ( .A(n2583), .Y(n8383) );
  DLY4X4 U9053 ( .A(n8387), .Y(n8386) );
  DLY4X4 U9054 ( .A(n3113), .Y(n8387) );
  AND2X1 U9055 ( .A(n2412), .B(N1658), .Y(n2291) );
  NAND3XL U9056 ( .A(n2587), .B(N1658), .C(n2586), .Y(n1461) );
  NOR3XL U9057 ( .A(n9512), .B(n9514), .C(n9511), .Y(n613) );
  NOR3XL U9058 ( .A(n9511), .B(n9512), .C(n9515), .Y(n1892) );
  NOR3XL U9059 ( .A(n9511), .B(n9514), .C(n9513), .Y(n1260) );
  INVX12 U9060 ( .A(n7241), .Y(IRB_A[2]) );
  INVX12 U9061 ( .A(n7242), .Y(IRB_A[3]) );
  INVX12 U9062 ( .A(n7243), .Y(IRB_A[4]) );
  INVX12 U9063 ( .A(n7244), .Y(IRB_A[5]) );
  INVX12 U9064 ( .A(n7246), .Y(IROM_A[5]) );
  NOR2BX2 U9065 ( .AN(n2536), .B(n9517), .Y(n667) );
  INVX3 U9066 ( .A(reset), .Y(n9669) );
  INVX3 U9067 ( .A(n2583), .Y(n8393) );
  MX4XL U9068 ( .A(n9173), .B(n9163), .C(n9168), .D(n9158), .S0(N1661), .S1(
        n8393), .Y(N7378) );
  MX4XL U9069 ( .A(n9193), .B(n9183), .C(n9188), .D(n9178), .S0(N1661), .S1(
        n8393), .Y(N7377) );
  MX4XL U9070 ( .A(n9213), .B(n9203), .C(n9208), .D(n9198), .S0(N1661), .S1(
        n8393), .Y(N7376) );
  MX4XL U9071 ( .A(n9233), .B(n9223), .C(n9228), .D(n9218), .S0(N1661), .S1(
        n8393), .Y(N7375) );
  MX4XL U9072 ( .A(n9253), .B(n9243), .C(n9248), .D(n9238), .S0(N1661), .S1(
        n8393), .Y(N7374) );
  MX4XL U9073 ( .A(n9273), .B(n9263), .C(n9268), .D(n9258), .S0(N1661), .S1(
        n8393), .Y(N7373) );
  OR2X1 U9079 ( .A(n2583), .B(n9339), .Y(n9831) );
  INVX12 U9080 ( .A(n9831), .Y(IROM_A[4]) );
  OR2X1 U9081 ( .A(n2586), .B(n9338), .Y(n9844) );
  INVX12 U9082 ( .A(n9844), .Y(IRB_A[1]) );
  OR2X1 U9083 ( .A(n2587), .B(n9338), .Y(n9845) );
  INVX12 U9084 ( .A(n9845), .Y(IRB_A[0]) );
  CLKBUFX3 U9085 ( .A(n2570), .Y(n9338) );
  BUFX12 U9086 ( .A(n9836), .Y(IRB_D[7]) );
  NOR2BX1 U9087 ( .AN(N7371), .B(n9338), .Y(n9836) );
  BUFX12 U9088 ( .A(n9837), .Y(IRB_D[6]) );
  NOR2BX1 U9089 ( .AN(N7372), .B(n9338), .Y(n9837) );
  BUFX12 U9090 ( .A(n9838), .Y(IRB_D[5]) );
  NOR2BX1 U9091 ( .AN(N7373), .B(n9338), .Y(n9838) );
  BUFX12 U9092 ( .A(n9839), .Y(IRB_D[4]) );
  NOR2BX1 U9093 ( .AN(N7374), .B(n9338), .Y(n9839) );
  BUFX12 U9094 ( .A(n9840), .Y(IRB_D[3]) );
  NOR2BX1 U9095 ( .AN(N7375), .B(n9338), .Y(n9840) );
  OR2X1 U9096 ( .A(n9339), .B(n2586), .Y(n9834) );
  INVX12 U9097 ( .A(n9834), .Y(IROM_A[1]) );
  CLKBUFX2 U9098 ( .A(n2563), .Y(n9339) );
  BUFX12 U9099 ( .A(n9841), .Y(IRB_D[2]) );
  NOR2BX1 U9100 ( .AN(N7376), .B(n9338), .Y(n9841) );
  OR2X1 U9101 ( .A(n9339), .B(n2585), .Y(n9833) );
  INVX12 U9102 ( .A(n9833), .Y(IROM_A[2]) );
  BUFX12 U9103 ( .A(n9846), .Y(busy) );
  BUFX12 U9104 ( .A(n9842), .Y(IRB_D[1]) );
  NOR2BX1 U9105 ( .AN(N7377), .B(n9338), .Y(n9842) );
  OR2X1 U9106 ( .A(n9339), .B(n2587), .Y(n9835) );
  INVX12 U9107 ( .A(n9835), .Y(IROM_A[0]) );
  BUFX12 U9108 ( .A(n9830), .Y(IROM_EN) );
  OR2X1 U9109 ( .A(n2584), .B(n9339), .Y(n9832) );
  INVX12 U9110 ( .A(n9832), .Y(IROM_A[3]) );
  BUFX12 U9111 ( .A(n9843), .Y(IRB_D[0]) );
  NOR2BX1 U9112 ( .AN(N7378), .B(n9338), .Y(n9843) );
  INVX16 U9113 ( .A(n2569), .Y(IRB_RW) );
  NAND2X1 U9114 ( .A(avg_reg[8]), .B(n9348), .Y(n280) );
  MX3XL U9115 ( .A(n8456), .B(n8903), .C(n8421), .S0(n8926), .S1(n8928), .Y(
        n8438) );
  OAI21XL U9116 ( .A0(n9666), .A1(n7225), .B0(n9625), .Y(n119) );
  CLKBUFX3 U9117 ( .A(n122), .Y(n9436) );
  OAI21XL U9118 ( .A0(n9664), .A1(n9621), .B0(n9618), .Y(n122) );
  CLKBUFX3 U9119 ( .A(n8931), .Y(n8936) );
  CLKBUFX3 U9120 ( .A(n8933), .Y(n8952) );
  CLKMX2X2 U9121 ( .A(n8510), .B(n8439), .S0(n8919), .Y(n8437) );
  CLKMX2X2 U9122 ( .A(n8438), .B(n8646), .S0(n8919), .Y(n8419) );
  MX3XL U9123 ( .A(n8457), .B(n8904), .C(n8422), .S0(n8926), .S1(n8928), .Y(
        n8439) );
  CLKMX2X2 U9124 ( .A(n8439), .B(n8659), .S0(n8919), .Y(n8420) );
  CLKBUFX3 U9125 ( .A(n9509), .Y(n8954) );
  MX4X1 U9126 ( .A(n8912), .B(n8422), .C(n8750), .D(n8746), .S0(n9127), .S1(
        n8929), .Y(n8418) );
  CLKMX2X2 U9127 ( .A(n8490), .B(n8438), .S0(n8919), .Y(n8436) );
  MXI3X1 U9128 ( .A(\buff[23][0] ), .B(\buff[27][0] ), .C(n8887), .S0(n8942), 
        .S1(n8958), .Y(n8491) );
  MXI3X1 U9129 ( .A(\buff[23][1] ), .B(\buff[27][1] ), .C(n8888), .S0(n8942), 
        .S1(n8958), .Y(n8511) );
  CLKBUFX3 U9130 ( .A(n273), .Y(n9632) );
  CLKBUFX3 U9131 ( .A(n287), .Y(n9623) );
  CLKBUFX3 U9132 ( .A(n273), .Y(n9630) );
  CLKBUFX3 U9133 ( .A(n287), .Y(n9621) );
  CLKBUFX3 U9134 ( .A(n273), .Y(n9631) );
  CLKBUFX3 U9135 ( .A(n287), .Y(n9622) );
  BUFX2 U9136 ( .A(n8932), .Y(n8933) );
  CLKBUFX3 U9137 ( .A(n266), .Y(n9638) );
  CLKBUFX3 U9138 ( .A(n266), .Y(n9637) );
  CLKINVX1 U9139 ( .A(n9514), .Y(n8920) );
  CLKBUFX3 U9140 ( .A(n9651), .Y(n9653) );
  CLKBUFX3 U9141 ( .A(n9645), .Y(n9647) );
  CLKBUFX3 U9142 ( .A(n9645), .Y(n9646) );
  CLKBUFX3 U9143 ( .A(n9657), .Y(n9659) );
  CLKBUFX3 U9144 ( .A(n9657), .Y(n9658) );
  CLKBUFX3 U9145 ( .A(n245), .Y(n9652) );
  INVX3 U9146 ( .A(n9386), .Y(n9781) );
  NAND3X2 U9147 ( .A(n9520), .B(n9376), .C(n2183), .Y(n2181) );
  NAND3X2 U9148 ( .A(n9524), .B(n9384), .C(n9376), .Y(n1862) );
  NAND3X2 U9149 ( .A(n9532), .B(n9414), .C(n9404), .Y(n910) );
  NAND3X2 U9150 ( .A(n9530), .B(n9404), .C(n9394), .Y(n1230) );
  NAND3X2 U9151 ( .A(n9526), .B(n9394), .C(n9384), .Y(n1547) );
  NAND3X2 U9152 ( .A(n9421), .B(n9424), .C(n9414), .Y(n582) );
  CLKINVX1 U9153 ( .A(n9510), .Y(n9138) );
  AOI22XL U9154 ( .A0(N7388), .A1(n9607), .B0(n8419), .B1(n9613), .Y(n624) );
  AO22XL U9155 ( .A0(n9433), .A1(n8419), .B0(n9434), .B1(N7388), .Y(n101) );
  AOI22X1 U9156 ( .A0(n9613), .A1(n8418), .B0(n9607), .B1(n8420), .Y(n8417) );
  CLKINVX1 U9157 ( .A(N7387), .Y(n9812) );
  CLKBUFX3 U9158 ( .A(n217), .Y(n9424) );
  CLKBUFX3 U9159 ( .A(n7245), .Y(n9522) );
  CLKINVX1 U9160 ( .A(N7386), .Y(n9811) );
  CLKINVX1 U9161 ( .A(N7385), .Y(n9810) );
  CLKINVX1 U9162 ( .A(N7384), .Y(n9809) );
  CLKINVX1 U9163 ( .A(N7383), .Y(n9808) );
  CLKINVX1 U9164 ( .A(N7382), .Y(n9807) );
  CLKINVX1 U9165 ( .A(N7381), .Y(n9806) );
  CLKINVX1 U9166 ( .A(N7380), .Y(n9805) );
  NAND3X2 U9167 ( .A(n9406), .B(n9407), .C(n9528), .Y(n1113) );
  NAND3X2 U9168 ( .A(n9377), .B(n9378), .C(n9518), .Y(n2099) );
  NAND3X2 U9169 ( .A(n9528), .B(n9398), .C(n9388), .Y(n1389) );
  NAND3X2 U9170 ( .A(n9518), .B(n9363), .C(n9364), .Y(n2382) );
  NAND3X2 U9171 ( .A(n2183), .B(n9358), .C(n9359), .Y(n2461) );
  NAND3X2 U9172 ( .A(n9414), .B(n9415), .C(n9405), .Y(n871) );
  NAND3X2 U9173 ( .A(n9395), .B(n9396), .C(n9781), .Y(n1469) );
  NAND3X2 U9174 ( .A(n9385), .B(n9781), .C(n9378), .Y(n1782) );
  NAND3X2 U9175 ( .A(n9404), .B(n9405), .C(n9395), .Y(n1191) );
  NAND3X2 U9176 ( .A(n9394), .B(n9395), .C(n9385), .Y(n1508) );
  NAND3X2 U9177 ( .A(n9384), .B(n9385), .C(n9377), .Y(n1823) );
  NAND3X2 U9178 ( .A(n9376), .B(n9377), .C(n9358), .Y(n2142) );
  NAND3X2 U9179 ( .A(n9781), .B(n9387), .C(n9379), .Y(n1743) );
  NAND3X2 U9180 ( .A(n9424), .B(n9425), .C(n9415), .Y(n542) );
  NAND3X2 U9181 ( .A(n9369), .B(n9371), .C(n9372), .Y(n2260) );
  NAND3X2 U9182 ( .A(n9366), .B(n9369), .C(n9370), .Y(n2302) );
  NAND3X2 U9183 ( .A(n9363), .B(n9366), .C(n9367), .Y(n2342) );
  NAND3X2 U9184 ( .A(n9419), .B(n9420), .C(n9410), .Y(n674) );
  NAND3X2 U9185 ( .A(n9418), .B(n9419), .C(n9409), .Y(n715) );
  NAND3X2 U9186 ( .A(n9417), .B(n9418), .C(n9408), .Y(n754) );
  NAND3X2 U9187 ( .A(n9416), .B(n9417), .C(n9407), .Y(n793) );
  NAND3X2 U9188 ( .A(n9415), .B(n9416), .C(n9406), .Y(n832) );
  NAND3X2 U9189 ( .A(n9409), .B(n9410), .C(n9400), .Y(n994) );
  NAND3X2 U9190 ( .A(n9408), .B(n9409), .C(n9399), .Y(n1035) );
  NAND3X2 U9191 ( .A(n9407), .B(n9408), .C(n9398), .Y(n1074) );
  NAND3X2 U9192 ( .A(n9405), .B(n9406), .C(n9396), .Y(n1152) );
  NAND3X2 U9193 ( .A(n9399), .B(n9400), .C(n9390), .Y(n1309) );
  NAND3X2 U9194 ( .A(n9398), .B(n9399), .C(n9389), .Y(n1350) );
  NAND3X2 U9195 ( .A(n9389), .B(n9390), .C(n9522), .Y(n1625) );
  NAND3X2 U9196 ( .A(n9380), .B(n9381), .C(n9369), .Y(n1982) );
  NAND3X2 U9197 ( .A(n9379), .B(n9380), .C(n9366), .Y(n2021) );
  NAND3X2 U9198 ( .A(n9378), .B(n9379), .C(n9363), .Y(n2060) );
  NAND3X2 U9199 ( .A(n9388), .B(n9389), .C(n9381), .Y(n1665) );
  NAND3X2 U9200 ( .A(n9387), .B(n9388), .C(n9380), .Y(n1704) );
  NAND3X2 U9201 ( .A(n9429), .B(n9430), .C(n9420), .Y(n309) );
  NAND3X2 U9202 ( .A(n9428), .B(n9429), .C(n9419), .Y(n382) );
  NAND3X2 U9203 ( .A(n9427), .B(n9428), .C(n9418), .Y(n422) );
  NAND3X2 U9204 ( .A(n9426), .B(n9427), .C(n9417), .Y(n462) );
  NAND3X2 U9205 ( .A(n9425), .B(n9426), .C(n9416), .Y(n502) );
  CLKBUFX2 U9206 ( .A(n9508), .Y(n9153) );
  BUFX2 U9207 ( .A(n9508), .Y(n8964) );
  CLKBUFX2 U9208 ( .A(n9508), .Y(n9152) );
  NAND2X1 U9209 ( .A(n2129), .B(n9349), .Y(n230) );
  NAND3X1 U9210 ( .A(N1656), .B(N1657), .C(n2291), .Y(n366) );
  CLKBUFX3 U9211 ( .A(n1577), .Y(n9344) );
  CLKBUFX3 U9212 ( .A(n613), .Y(n9411) );
  CLKBUFX3 U9213 ( .A(n940), .Y(n9401) );
  CLKBUFX3 U9214 ( .A(n151), .Y(n9429) );
  CLKBUFX3 U9215 ( .A(n165), .Y(n9428) );
  CLKBUFX3 U9216 ( .A(n178), .Y(n9427) );
  CLKBUFX3 U9217 ( .A(n191), .Y(n9426) );
  CLKBUFX3 U9218 ( .A(n204), .Y(n9425) );
  AOI221XL U9219 ( .A0(n8373), .A1(n2557), .B0(n9516), .B1(n2552), .C0(n2549), 
        .Y(n2551) );
  BUFX4 U9220 ( .A(n312), .Y(n9420) );
  MX4XL U9221 ( .A(\buff[8][2] ), .B(\buff[12][2] ), .C(\buff[10][2] ), .D(
        \buff[14][2] ), .S0(n8951), .S1(n8416), .Y(n8519) );
  MX4XL U9222 ( .A(\buff[40][2] ), .B(\buff[44][2] ), .C(\buff[42][2] ), .D(
        \buff[46][2] ), .S0(n8951), .S1(n9145), .Y(n8518) );
  MX4XL U9223 ( .A(\buff[8][3] ), .B(\buff[12][3] ), .C(\buff[10][3] ), .D(
        \buff[14][3] ), .S0(n8951), .S1(n9144), .Y(n8539) );
  MX4XL U9224 ( .A(\buff[40][3] ), .B(\buff[44][3] ), .C(\buff[42][3] ), .D(
        \buff[46][3] ), .S0(n8951), .S1(n9143), .Y(n8538) );
  MXI2XL U9225 ( .A(\buff[25][2] ), .B(\buff[29][2] ), .S0(n8431), .Y(n8670)
         );
  MXI2XL U9226 ( .A(\buff[1][0] ), .B(\buff[5][0] ), .S0(n8947), .Y(n8487) );
  MXI2XL U9227 ( .A(\buff[1][1] ), .B(\buff[5][1] ), .S0(n8947), .Y(n8507) );
  MXI2XL U9228 ( .A(\buff[1][2] ), .B(\buff[5][2] ), .S0(n8431), .Y(n8527) );
  MXI2XL U9229 ( .A(\buff[49][0] ), .B(\buff[53][0] ), .S0(n8947), .Y(n8481)
         );
  MXI2XL U9230 ( .A(\buff[49][1] ), .B(\buff[53][1] ), .S0(n8947), .Y(n8501)
         );
  MXI2XL U9231 ( .A(\buff[33][1] ), .B(\buff[37][1] ), .S0(n8947), .Y(n8505)
         );
  MXI2XL U9232 ( .A(\buff[33][0] ), .B(\buff[37][0] ), .S0(n8947), .Y(n8485)
         );
  MXI2XL U9233 ( .A(\buff[33][2] ), .B(\buff[37][2] ), .S0(n8431), .Y(n8525)
         );
  MXI2XL U9234 ( .A(\buff[49][2] ), .B(\buff[53][2] ), .S0(n8431), .Y(n8521)
         );
  MXI2XL U9235 ( .A(\buff[17][0] ), .B(\buff[21][0] ), .S0(n8947), .Y(n8483)
         );
  MXI2XL U9236 ( .A(\buff[17][1] ), .B(\buff[21][1] ), .S0(n8947), .Y(n8503)
         );
  MXI2XL U9237 ( .A(\buff[17][2] ), .B(\buff[21][2] ), .S0(n8431), .Y(n8523)
         );
  MXI2XL U9238 ( .A(\buff[41][0] ), .B(\buff[45][0] ), .S0(n8947), .Y(n8488)
         );
  MXI2XL U9239 ( .A(\buff[41][1] ), .B(\buff[45][1] ), .S0(n8947), .Y(n8508)
         );
  MXI2XL U9240 ( .A(\buff[9][0] ), .B(\buff[13][0] ), .S0(n8947), .Y(n8489) );
  MXI2XL U9241 ( .A(\buff[9][1] ), .B(\buff[13][1] ), .S0(n8947), .Y(n8509) );
  MX4XL U9242 ( .A(\buff[56][2] ), .B(\buff[60][2] ), .C(\buff[58][2] ), .D(
        \buff[62][2] ), .S0(n8948), .S1(n8959), .Y(n8752) );
  MX4XL U9243 ( .A(\buff[55][1] ), .B(\buff[59][1] ), .C(\buff[57][1] ), .D(
        \buff[61][1] ), .S0(n8949), .S1(n8959), .Y(n8749) );
  MX4XL U9244 ( .A(\buff[55][0] ), .B(\buff[59][0] ), .C(\buff[57][0] ), .D(
        \buff[61][0] ), .S0(n8949), .S1(n8959), .Y(n8742) );
  INVX1 U9245 ( .A(n8644), .Y(n8887) );
  INVX1 U9246 ( .A(n8657), .Y(n8888) );
  MX4X1 U9247 ( .A(n8477), .B(n8475), .C(n8476), .D(n8474), .S0(n8926), .S1(
        n8922), .Y(n8421) );
  MX4X1 U9248 ( .A(n8497), .B(n8495), .C(n8496), .D(n8494), .S0(n8926), .S1(
        n8922), .Y(n8422) );
  MX4X1 U9249 ( .A(n8517), .B(n8515), .C(n8516), .D(n8514), .S0(n8926), .S1(
        n8922), .Y(n8423) );
  MX4X1 U9250 ( .A(n8537), .B(n8535), .C(n8536), .D(n8534), .S0(n8927), .S1(
        n8922), .Y(n8424) );
  MXI4XL U9251 ( .A(n8487), .B(n8638), .C(n8485), .D(n8639), .S0(n8961), .S1(
        n8923), .Y(n8637) );
  MXI4XL U9252 ( .A(n8483), .B(n8635), .C(n8481), .D(n8636), .S0(n8961), .S1(
        n8922), .Y(n8634) );
  MXI4XL U9253 ( .A(n8503), .B(n8648), .C(n8501), .D(n8649), .S0(n8962), .S1(
        n8921), .Y(n8647) );
  MXI4XL U9254 ( .A(n8507), .B(n8651), .C(n8505), .D(n8652), .S0(n8961), .S1(
        n8921), .Y(n8650) );
  MX4XL U9255 ( .A(\buff[0][1] ), .B(\buff[4][1] ), .C(\buff[2][1] ), .D(
        \buff[6][1] ), .S0(n8952), .S1(n8416), .Y(n8497) );
  MX4XL U9256 ( .A(\buff[0][2] ), .B(\buff[4][2] ), .C(\buff[2][2] ), .D(
        \buff[6][2] ), .S0(n8951), .S1(n9144), .Y(n8517) );
  MX4XL U9257 ( .A(\buff[0][3] ), .B(\buff[4][3] ), .C(\buff[2][3] ), .D(
        \buff[6][3] ), .S0(n8951), .S1(n9142), .Y(n8537) );
  MX4XL U9258 ( .A(\buff[16][1] ), .B(\buff[20][1] ), .C(\buff[18][1] ), .D(
        \buff[22][1] ), .S0(n8952), .S1(n8416), .Y(n8495) );
  MX4XL U9259 ( .A(\buff[16][2] ), .B(\buff[20][2] ), .C(\buff[18][2] ), .D(
        \buff[22][2] ), .S0(n8951), .S1(n9144), .Y(n8515) );
  MX4XL U9260 ( .A(\buff[16][3] ), .B(\buff[20][3] ), .C(\buff[18][3] ), .D(
        \buff[22][3] ), .S0(n8951), .S1(n9143), .Y(n8535) );
  MX4XL U9261 ( .A(\buff[8][4] ), .B(\buff[12][4] ), .C(\buff[10][4] ), .D(
        \buff[14][4] ), .S0(n8950), .S1(n9142), .Y(n8559) );
  MX4XL U9262 ( .A(\buff[40][4] ), .B(\buff[44][4] ), .C(\buff[42][4] ), .D(
        \buff[46][4] ), .S0(n8950), .S1(n9148), .Y(n8558) );
  MX4XL U9263 ( .A(\buff[8][5] ), .B(\buff[12][5] ), .C(\buff[10][5] ), .D(
        \buff[14][5] ), .S0(n8950), .S1(n9150), .Y(n8579) );
  MX4XL U9264 ( .A(\buff[40][5] ), .B(\buff[44][5] ), .C(\buff[42][5] ), .D(
        \buff[46][5] ), .S0(n8950), .S1(n9150), .Y(n8578) );
  MX4X1 U9265 ( .A(n8577), .B(n8575), .C(n8576), .D(n8574), .S0(n8926), .S1(
        n8923), .Y(n8425) );
  MX4X1 U9266 ( .A(n8557), .B(n8555), .C(n8556), .D(n8554), .S0(n8927), .S1(
        n8922), .Y(n8426) );
  MX4XL U9267 ( .A(\buff[0][4] ), .B(\buff[4][4] ), .C(\buff[2][4] ), .D(
        \buff[6][4] ), .S0(n8950), .S1(n9142), .Y(n8557) );
  MX4XL U9268 ( .A(\buff[0][5] ), .B(\buff[4][5] ), .C(\buff[2][5] ), .D(
        \buff[6][5] ), .S0(n8950), .S1(n9151), .Y(n8577) );
  MX4XL U9269 ( .A(\buff[16][4] ), .B(\buff[20][4] ), .C(\buff[18][4] ), .D(
        \buff[22][4] ), .S0(n8951), .S1(n9142), .Y(n8555) );
  MX4XL U9270 ( .A(\buff[16][5] ), .B(\buff[20][5] ), .C(\buff[18][5] ), .D(
        \buff[22][5] ), .S0(n8950), .S1(n9151), .Y(n8575) );
  MX4XL U9271 ( .A(\buff[8][6] ), .B(\buff[12][6] ), .C(\buff[10][6] ), .D(
        \buff[14][6] ), .S0(n8949), .S1(n9146), .Y(n8599) );
  MX4XL U9272 ( .A(\buff[40][6] ), .B(\buff[44][6] ), .C(\buff[42][6] ), .D(
        \buff[46][6] ), .S0(n8949), .S1(n8958), .Y(n8598) );
  MX4XL U9273 ( .A(\buff[8][7] ), .B(\buff[12][7] ), .C(\buff[10][7] ), .D(
        \buff[14][7] ), .S0(n8949), .S1(n9145), .Y(n8619) );
  AOI211XL U9274 ( .A0(n233), .A1(n8436), .B0(n234), .C0(n9450), .Y(n232) );
  INVXL U9275 ( .A(n8436), .Y(n9804) );
  AOI211XL U9276 ( .A0(n233), .A1(n8437), .B0(n244), .C0(n9448), .Y(n243) );
  INVXL U9277 ( .A(n8437), .Y(n9803) );
  MX4XL U9278 ( .A(\buff[56][5] ), .B(\buff[60][5] ), .C(\buff[58][5] ), .D(
        \buff[62][5] ), .S0(n8948), .S1(n9145), .Y(n8773) );
  MX4X1 U9279 ( .A(n8597), .B(n8595), .C(n8596), .D(n8594), .S0(n8927), .S1(
        n8923), .Y(n8427) );
  MX4X1 U9280 ( .A(n8617), .B(n8615), .C(n8616), .D(n8614), .S0(n8927), .S1(
        n8923), .Y(n8428) );
  MX4XL U9281 ( .A(\buff[0][6] ), .B(\buff[4][6] ), .C(\buff[2][6] ), .D(
        \buff[6][6] ), .S0(n8949), .S1(n8956), .Y(n8597) );
  MX4XL U9282 ( .A(\buff[0][7] ), .B(\buff[4][7] ), .C(\buff[2][7] ), .D(
        \buff[6][7] ), .S0(n8949), .S1(n9145), .Y(n8617) );
  MX4XL U9283 ( .A(\buff[16][6] ), .B(\buff[20][6] ), .C(\buff[18][6] ), .D(
        \buff[22][6] ), .S0(n8950), .S1(n8963), .Y(n8595) );
  MX4XL U9284 ( .A(\buff[16][7] ), .B(\buff[20][7] ), .C(\buff[18][7] ), .D(
        \buff[22][7] ), .S0(n8949), .S1(n9143), .Y(n8615) );
  NOR2X2 U9285 ( .A(n9741), .B(reset), .Y(n2129) );
  NAND3X1 U9286 ( .A(n2586), .B(n2587), .C(n2132), .Y(n299) );
  CLKBUFX3 U9287 ( .A(n1421), .Y(n9397) );
  CLKBUFX3 U9288 ( .A(n2415), .Y(n9360) );
  NOR2X1 U9289 ( .A(n9666), .B(n8372), .Y(n985) );
  NAND3X1 U9290 ( .A(n9744), .B(n2581), .C(N1677), .Y(n982) );
  CLKBUFX3 U9291 ( .A(n375), .Y(n9341) );
  NOR3XL U9292 ( .A(n2576), .B(n2575), .C(n9516), .Y(n375) );
  NOR3X1 U9293 ( .A(n9738), .B(n2590), .C(n9747), .Y(n2541) );
  NOR3X1 U9294 ( .A(n9738), .B(n2589), .C(n9748), .Y(n2552) );
  CLKBUFX3 U9295 ( .A(n415), .Y(n9368) );
  NOR3XL U9296 ( .A(n2576), .B(n2575), .C(n9517), .Y(n415) );
  CLKBUFX3 U9297 ( .A(n455), .Y(n9365) );
  NOR3XL U9298 ( .A(n9516), .B(n2575), .C(n9508), .Y(n455) );
  CLKBUFX3 U9299 ( .A(n575), .Y(n9357) );
  NOR3XL U9300 ( .A(n9517), .B(n2576), .C(n9509), .Y(n575) );
  CLKBUFX3 U9301 ( .A(n495), .Y(n9362) );
  NOR3XL U9302 ( .A(n9517), .B(n2575), .C(n9508), .Y(n495) );
  CLKBUFX3 U9303 ( .A(n535), .Y(n9342) );
  NOR3XL U9304 ( .A(n9516), .B(n2576), .C(n9509), .Y(n535) );
  NOR4X1 U9305 ( .A(n9339), .B(n9340), .C(n981), .D(n2581), .Y(n96) );
  NOR3BX1 U9306 ( .AN(n2581), .B(n1975), .C(n159), .Y(n91) );
  OAI2BB2XL U9307 ( .B0(n9457), .B1(n140), .A0N(n7318), .A1N(n9457), .Y(n2608)
         );
  AND2X2 U9308 ( .A(n9796), .B(n141), .Y(n8429) );
  AND2X2 U9309 ( .A(n9437), .B(n9430), .Y(n8430) );
  NOR3XL U9310 ( .A(n8429), .B(n8430), .C(n9438), .Y(n140) );
  CLKBUFX2 U9311 ( .A(n9509), .Y(n9141) );
  CLKBUFX3 U9312 ( .A(n9126), .Y(n9135) );
  CLKBUFX3 U9313 ( .A(n9126), .Y(n9134) );
  CLKBUFX3 U9314 ( .A(n9127), .Y(n9133) );
  CLKBUFX3 U9315 ( .A(n9128), .Y(n9132) );
  CLKBUFX3 U9316 ( .A(n9129), .Y(n9131) );
  CLKBUFX3 U9317 ( .A(n9131), .Y(n9130) );
  CLKBUFX3 U9318 ( .A(n9481), .Y(n9482) );
  CLKBUFX3 U9319 ( .A(n9732), .Y(n9478) );
  CLKBUFX3 U9320 ( .A(n9731), .Y(n9475) );
  CLKBUFX3 U9321 ( .A(n9730), .Y(n9472) );
  CLKBUFX3 U9322 ( .A(n9729), .Y(n9469) );
  CLKBUFX3 U9323 ( .A(n9728), .Y(n9466) );
  CLKBUFX3 U9324 ( .A(n9727), .Y(n9463) );
  CLKBUFX3 U9325 ( .A(n9726), .Y(n9460) );
  CLKBUFX3 U9326 ( .A(n9481), .Y(n9483) );
  CLKBUFX3 U9327 ( .A(n9732), .Y(n9479) );
  CLKBUFX3 U9328 ( .A(n9731), .Y(n9476) );
  CLKBUFX3 U9329 ( .A(n9730), .Y(n9473) );
  CLKBUFX3 U9330 ( .A(n9729), .Y(n9470) );
  CLKBUFX3 U9331 ( .A(n9728), .Y(n9467) );
  CLKBUFX3 U9332 ( .A(n9727), .Y(n9464) );
  CLKBUFX3 U9333 ( .A(n9726), .Y(n9461) );
  CLKBUFX3 U9334 ( .A(n9732), .Y(n9480) );
  CLKBUFX3 U9335 ( .A(n9731), .Y(n9477) );
  CLKBUFX3 U9336 ( .A(n9730), .Y(n9474) );
  CLKBUFX3 U9337 ( .A(n9729), .Y(n9471) );
  CLKBUFX3 U9338 ( .A(n9728), .Y(n9468) );
  CLKBUFX3 U9339 ( .A(n9727), .Y(n9465) );
  CLKBUFX3 U9340 ( .A(n9726), .Y(n9462) );
  OAI21XL U9341 ( .A0(n9576), .A1(n2181), .B0(n7226), .Y(n2195) );
  OAI21XL U9342 ( .A0(n9567), .A1(n2181), .B0(n9636), .Y(n2199) );
  OAI21XL U9343 ( .A0(n9560), .A1(n2181), .B0(n9630), .Y(n2203) );
  OAI21XL U9344 ( .A0(n9550), .A1(n2181), .B0(n7225), .Y(n2207) );
  OAI21XL U9345 ( .A0(n9540), .A1(n2181), .B0(n9622), .Y(n2213) );
  OAI21XL U9346 ( .A0(n9578), .A1(n582), .B0(n7226), .Y(n596) );
  OAI21XL U9347 ( .A0(n9569), .A1(n582), .B0(n9638), .Y(n600) );
  OAI21XL U9348 ( .A0(n9560), .A1(n582), .B0(n9632), .Y(n604) );
  OAI21XL U9349 ( .A0(n9550), .A1(n582), .B0(n7225), .Y(n608) );
  OAI21XL U9350 ( .A0(n9542), .A1(n582), .B0(n9623), .Y(n616) );
  OAI21XL U9351 ( .A0(n9577), .A1(n910), .B0(n7226), .Y(n924) );
  OAI21XL U9352 ( .A0(n9568), .A1(n910), .B0(n9637), .Y(n928) );
  OAI21XL U9353 ( .A0(n9559), .A1(n910), .B0(n9631), .Y(n932) );
  OAI21XL U9354 ( .A0(n9549), .A1(n910), .B0(n7225), .Y(n936) );
  OAI21XL U9355 ( .A0(n9540), .A1(n910), .B0(n9622), .Y(n942) );
  OAI21XL U9356 ( .A0(n9577), .A1(n1230), .B0(n7226), .Y(n1244) );
  OAI21XL U9357 ( .A0(n9568), .A1(n1230), .B0(n9637), .Y(n1248) );
  OAI21XL U9358 ( .A0(n9559), .A1(n1230), .B0(n9631), .Y(n1252) );
  OAI21XL U9359 ( .A0(n9549), .A1(n1230), .B0(n7225), .Y(n1256) );
  OAI21XL U9360 ( .A0(n9540), .A1(n1230), .B0(n9622), .Y(n1262) );
  OAI21XL U9361 ( .A0(n9578), .A1(n1547), .B0(n7226), .Y(n1561) );
  OAI21XL U9362 ( .A0(n9568), .A1(n1547), .B0(n9637), .Y(n1565) );
  OAI21XL U9363 ( .A0(n9558), .A1(n1547), .B0(n9630), .Y(n1569) );
  OAI21XL U9364 ( .A0(n9551), .A1(n1547), .B0(n7225), .Y(n1573) );
  OAI21XL U9365 ( .A0(n9541), .A1(n1547), .B0(n9621), .Y(n1579) );
  OAI21XL U9366 ( .A0(n9576), .A1(n1862), .B0(n7226), .Y(n1876) );
  OAI21XL U9367 ( .A0(n9567), .A1(n1862), .B0(n9637), .Y(n1880) );
  OAI21XL U9368 ( .A0(n9559), .A1(n1862), .B0(n9630), .Y(n1884) );
  OAI21XL U9369 ( .A0(n9551), .A1(n1862), .B0(n7225), .Y(n1888) );
  OAI21XL U9370 ( .A0(n9540), .A1(n1862), .B0(n9621), .Y(n1894) );
  CLKBUFX3 U9371 ( .A(n8934), .Y(n8951) );
  CLKBUFX3 U9372 ( .A(n8935), .Y(n8949) );
  CLKBUFX3 U9373 ( .A(n8936), .Y(n8947) );
  CLKBUFX3 U9374 ( .A(n8938), .Y(n8945) );
  CLKBUFX3 U9375 ( .A(n8925), .Y(n8926) );
  CLKBUFX3 U9376 ( .A(n9125), .Y(n9126) );
  OAI21XL U9377 ( .A0(n9603), .A1(n2181), .B0(n9657), .Y(n2180) );
  OAI21XL U9378 ( .A0(n9595), .A1(n2181), .B0(n9651), .Y(n2187) );
  OAI21XL U9379 ( .A0(n9587), .A1(n2181), .B0(n252), .Y(n2191) );
  OAI21XL U9380 ( .A0(n9604), .A1(n582), .B0(n9659), .Y(n581) );
  OAI21XL U9381 ( .A0(n9596), .A1(n582), .B0(n9653), .Y(n588) );
  OAI21XL U9382 ( .A0(n9587), .A1(n582), .B0(n9647), .Y(n592) );
  OAI21XL U9383 ( .A0(n9605), .A1(n910), .B0(n9658), .Y(n909) );
  OAI21XL U9384 ( .A0(n9595), .A1(n910), .B0(n9652), .Y(n916) );
  OAI21XL U9385 ( .A0(n9586), .A1(n910), .B0(n9646), .Y(n920) );
  OAI21XL U9386 ( .A0(n9605), .A1(n1230), .B0(n9658), .Y(n1229) );
  OAI21XL U9387 ( .A0(n9595), .A1(n1230), .B0(n9652), .Y(n1236) );
  OAI21XL U9388 ( .A0(n9586), .A1(n1230), .B0(n252), .Y(n1240) );
  OAI21XL U9389 ( .A0(n9605), .A1(n1547), .B0(n9658), .Y(n1546) );
  OAI21XL U9390 ( .A0(n9595), .A1(n1547), .B0(n9652), .Y(n1553) );
  OAI21XL U9391 ( .A0(n9585), .A1(n1547), .B0(n9646), .Y(n1557) );
  OAI21XL U9392 ( .A0(n9603), .A1(n1862), .B0(n9658), .Y(n1861) );
  OAI21XL U9393 ( .A0(n9594), .A1(n1862), .B0(n9652), .Y(n1868) );
  OAI21XL U9394 ( .A0(n9586), .A1(n1862), .B0(n9646), .Y(n1872) );
  CLKBUFX3 U9395 ( .A(n8934), .Y(n8950) );
  CLKBUFX3 U9396 ( .A(n8935), .Y(n8948) );
  CLKBUFX3 U9397 ( .A(n8937), .Y(n8946) );
  CLKBUFX3 U9398 ( .A(n8924), .Y(n8927) );
  BUFX4 U9399 ( .A(n8920), .Y(n8922) );
  CLKBUFX3 U9400 ( .A(n8920), .Y(n8923) );
  CLKBUFX3 U9401 ( .A(n8920), .Y(n8921) );
  CLKBUFX3 U9402 ( .A(n9125), .Y(n9127) );
  CLKBUFX3 U9403 ( .A(n9125), .Y(n9128) );
  CLKBUFX3 U9404 ( .A(n9128), .Y(n9129) );
  CLKBUFX3 U9405 ( .A(n308), .Y(n9604) );
  CLKBUFX3 U9406 ( .A(n9594), .Y(n9596) );
  CLKBUFX3 U9407 ( .A(n7240), .Y(n9587) );
  CLKBUFX3 U9408 ( .A(n7239), .Y(n9578) );
  CLKBUFX3 U9409 ( .A(n7237), .Y(n9569) );
  CLKBUFX3 U9410 ( .A(n351), .Y(n9560) );
  CLKBUFX3 U9411 ( .A(n7238), .Y(n9550) );
  CLKBUFX3 U9412 ( .A(n7232), .Y(n9542) );
  CLKBUFX3 U9413 ( .A(n313), .Y(n9598) );
  CLKBUFX3 U9414 ( .A(n321), .Y(n9589) );
  CLKBUFX3 U9415 ( .A(n329), .Y(n9580) );
  CLKBUFX3 U9416 ( .A(n337), .Y(n9571) );
  CLKBUFX3 U9417 ( .A(n353), .Y(n9553) );
  CLKBUFX3 U9418 ( .A(n361), .Y(n9544) );
  CLKBUFX3 U9419 ( .A(n374), .Y(n9535) );
  CLKBUFX3 U9420 ( .A(n313), .Y(n9599) );
  CLKBUFX3 U9421 ( .A(n9579), .Y(n9581) );
  CLKBUFX3 U9422 ( .A(n9570), .Y(n9572) );
  CLKBUFX3 U9423 ( .A(n9561), .Y(n9563) );
  CLKBUFX3 U9424 ( .A(n353), .Y(n9554) );
  CLKBUFX3 U9425 ( .A(n361), .Y(n9545) );
  CLKBUFX3 U9426 ( .A(n374), .Y(n9536) );
  CLKBUFX3 U9427 ( .A(n313), .Y(n9597) );
  CLKBUFX3 U9428 ( .A(n321), .Y(n9588) );
  CLKBUFX3 U9429 ( .A(n329), .Y(n9579) );
  CLKBUFX3 U9430 ( .A(n337), .Y(n9570) );
  CLKBUFX3 U9431 ( .A(n345), .Y(n9562) );
  CLKBUFX3 U9432 ( .A(n353), .Y(n9552) );
  CLKBUFX3 U9433 ( .A(n361), .Y(n9543) );
  CLKBUFX3 U9434 ( .A(n374), .Y(n9534) );
  CLKBUFX3 U9435 ( .A(n9586), .Y(n9585) );
  CLKBUFX3 U9436 ( .A(n351), .Y(n9558) );
  CLKBUFX3 U9437 ( .A(n7232), .Y(n9541) );
  CLKBUFX3 U9438 ( .A(n9594), .Y(n9595) );
  CLKBUFX3 U9439 ( .A(n7240), .Y(n9586) );
  CLKBUFX3 U9440 ( .A(n7239), .Y(n9577) );
  CLKBUFX3 U9441 ( .A(n7237), .Y(n9568) );
  CLKBUFX3 U9442 ( .A(n351), .Y(n9559) );
  CLKBUFX3 U9443 ( .A(n7238), .Y(n9549) );
  CLKBUFX3 U9444 ( .A(n9605), .Y(n9603) );
  CLKBUFX3 U9445 ( .A(n9577), .Y(n9576) );
  CLKBUFX3 U9446 ( .A(n7232), .Y(n9540) );
  CLKBUFX3 U9447 ( .A(n9591), .Y(n9592) );
  CLKBUFX3 U9448 ( .A(n9582), .Y(n9583) );
  CLKBUFX3 U9449 ( .A(n9573), .Y(n9574) );
  CLKBUFX3 U9450 ( .A(n360), .Y(n9546) );
  CLKBUFX3 U9451 ( .A(n373), .Y(n9537) );
  CLKBUFX3 U9452 ( .A(n310), .Y(n9600) );
  CLKBUFX3 U9453 ( .A(n9591), .Y(n9593) );
  CLKBUFX3 U9454 ( .A(n9582), .Y(n9584) );
  CLKBUFX3 U9455 ( .A(n9573), .Y(n9575) );
  CLKBUFX3 U9456 ( .A(n9564), .Y(n9565) );
  CLKBUFX3 U9457 ( .A(n352), .Y(n9555) );
  CLKBUFX3 U9458 ( .A(n360), .Y(n9547) );
  CLKBUFX3 U9459 ( .A(n373), .Y(n9538) );
  CLKBUFX3 U9460 ( .A(n310), .Y(n9602) );
  CLKBUFX3 U9461 ( .A(n352), .Y(n9557) );
  CLKBUFX3 U9462 ( .A(n360), .Y(n9548) );
  CLKBUFX3 U9463 ( .A(n373), .Y(n9539) );
  CLKBUFX3 U9464 ( .A(n310), .Y(n9601) );
  CLKBUFX3 U9465 ( .A(n9564), .Y(n9566) );
  CLKBUFX3 U9466 ( .A(n352), .Y(n9556) );
  CLKBUFX3 U9467 ( .A(n9733), .Y(n9481) );
  CLKBUFX3 U9468 ( .A(n9588), .Y(n9590) );
  CLKBUFX3 U9469 ( .A(n9316), .Y(n9318) );
  CLKBUFX3 U9470 ( .A(n9316), .Y(n9319) );
  CLKBUFX3 U9471 ( .A(n9315), .Y(n9321) );
  CLKBUFX3 U9472 ( .A(n9316), .Y(n9320) );
  CLKBUFX3 U9473 ( .A(n9315), .Y(n9322) );
  CLKBUFX3 U9474 ( .A(n9314), .Y(n9323) );
  CLKBUFX3 U9475 ( .A(n9314), .Y(n9324) );
  CLKBUFX3 U9476 ( .A(n9315), .Y(n9317) );
  OAI221XL U9477 ( .A0(n1428), .A1(n9496), .B0(n9578), .B1(n1429), .C0(n7226), 
        .Y(n1440) );
  OAI221XL U9478 ( .A0(n1428), .A1(n9808), .B0(n9569), .B1(n1429), .C0(n9638), 
        .Y(n1444) );
  OAI221XL U9479 ( .A0(n1428), .A1(n9490), .B0(n9560), .B1(n1429), .C0(n9632), 
        .Y(n1448) );
  OAI221XL U9480 ( .A0(n1428), .A1(n9487), .B0(n9550), .B1(n1429), .C0(n7225), 
        .Y(n1452) );
  OAI221XL U9481 ( .A0(n1428), .A1(n9484), .B0(n9542), .B1(n1429), .C0(n9623), 
        .Y(n1456) );
  OAI221XL U9482 ( .A0(n1941), .A1(n9809), .B0(n9578), .B1(n1942), .C0(n7226), 
        .Y(n1953) );
  OAI221XL U9483 ( .A0(n1941), .A1(n9808), .B0(n9569), .B1(n1942), .C0(n9638), 
        .Y(n1957) );
  OAI221XL U9484 ( .A0(n1941), .A1(n9490), .B0(n9560), .B1(n1942), .C0(n9632), 
        .Y(n1961) );
  OAI221XL U9485 ( .A0(n1941), .A1(n9487), .B0(n9550), .B1(n1942), .C0(n7225), 
        .Y(n1965) );
  OAI221XL U9486 ( .A0(n1941), .A1(n9484), .B0(n9542), .B1(n1942), .C0(n9623), 
        .Y(n1969) );
  OAI221XL U9487 ( .A0(n2422), .A1(n9493), .B0(n9567), .B1(n2423), .C0(n9637), 
        .Y(n2438) );
  OAI221XL U9488 ( .A0(n2422), .A1(n9490), .B0(n9558), .B1(n2423), .C0(n9630), 
        .Y(n2442) );
  OAI221XL U9489 ( .A0(n2422), .A1(n9487), .B0(n9551), .B1(n2423), .C0(n7225), 
        .Y(n2446) );
  OAI221XL U9490 ( .A0(n2422), .A1(n9484), .B0(n7232), .B1(n2423), .C0(n9621), 
        .Y(n2450) );
  OAI221XL U9491 ( .A0(n1902), .A1(n9495), .B0(n9567), .B1(n1903), .C0(n9637), 
        .Y(n1918) );
  OAI221XL U9492 ( .A0(n1902), .A1(n9490), .B0(n9558), .B1(n1903), .C0(n9631), 
        .Y(n1922) );
  OAI221XL U9493 ( .A0(n1902), .A1(n9487), .B0(n9551), .B1(n1903), .C0(n7225), 
        .Y(n1926) );
  OAI221XL U9494 ( .A0(n1902), .A1(n9484), .B0(n7232), .B1(n1903), .C0(n9622), 
        .Y(n1930) );
  OAI221XL U9495 ( .A0(n626), .A1(n9498), .B0(n9578), .B1(n9422), .C0(n7226), 
        .Y(n640) );
  OAI221XL U9496 ( .A0(n626), .A1(n9495), .B0(n9567), .B1(n9422), .C0(n9638), 
        .Y(n645) );
  OAI221XL U9497 ( .A0(n626), .A1(n9490), .B0(n9559), .B1(n9422), .C0(n9632), 
        .Y(n650) );
  OAI221XL U9498 ( .A0(n626), .A1(n9487), .B0(n9551), .B1(n9422), .C0(n7225), 
        .Y(n655) );
  OAI221XL U9499 ( .A0(n626), .A1(n9484), .B0(n9542), .B1(n9422), .C0(n9623), 
        .Y(n660) );
  OAI221XL U9500 ( .A0(n950), .A1(n9498), .B0(n9578), .B1(n9412), .C0(n7226), 
        .Y(n962) );
  OAI221XL U9501 ( .A0(n950), .A1(n9494), .B0(n9569), .B1(n9412), .C0(n9638), 
        .Y(n966) );
  OAI221XL U9502 ( .A0(n950), .A1(n9490), .B0(n9560), .B1(n9412), .C0(n9632), 
        .Y(n970) );
  OAI221XL U9503 ( .A0(n950), .A1(n9487), .B0(n9550), .B1(n9412), .C0(n7225), 
        .Y(n974) );
  OAI221XL U9504 ( .A0(n950), .A1(n9484), .B0(n9542), .B1(n9412), .C0(n9623), 
        .Y(n978) );
  OAI221XL U9505 ( .A0(n1270), .A1(n9496), .B0(n9578), .B1(n9402), .C0(n7226), 
        .Y(n1282) );
  OAI221XL U9506 ( .A0(n1270), .A1(n9494), .B0(n9569), .B1(n9402), .C0(n9638), 
        .Y(n1286) );
  OAI221XL U9507 ( .A0(n1270), .A1(n9490), .B0(n9560), .B1(n9402), .C0(n9632), 
        .Y(n1290) );
  OAI221XL U9508 ( .A0(n1270), .A1(n9487), .B0(n9550), .B1(n9402), .C0(n7225), 
        .Y(n1294) );
  OAI221XL U9509 ( .A0(n1270), .A1(n9484), .B0(n9542), .B1(n9402), .C0(n9623), 
        .Y(n1298) );
  OAI221XL U9510 ( .A0(n1587), .A1(n9809), .B0(n9578), .B1(n9392), .C0(n7226), 
        .Y(n1599) );
  OAI221XL U9511 ( .A0(n1587), .A1(n9808), .B0(n9569), .B1(n9392), .C0(n9638), 
        .Y(n1603) );
  OAI221XL U9512 ( .A0(n1587), .A1(n9490), .B0(n9560), .B1(n9392), .C0(n9632), 
        .Y(n1607) );
  OAI221XL U9513 ( .A0(n1587), .A1(n9487), .B0(n9550), .B1(n9392), .C0(n7225), 
        .Y(n1611) );
  OAI221XL U9514 ( .A0(n1587), .A1(n9484), .B0(n9542), .B1(n9392), .C0(n9623), 
        .Y(n1615) );
  OAI221XL U9515 ( .A0(n2221), .A1(n9809), .B0(n9577), .B1(n9374), .C0(n7226), 
        .Y(n2233) );
  OAI221XL U9516 ( .A0(n2221), .A1(n9808), .B0(n9567), .B1(n9374), .C0(n9638), 
        .Y(n2237) );
  OAI221XL U9517 ( .A0(n2221), .A1(n9490), .B0(n9559), .B1(n9374), .C0(n9632), 
        .Y(n2241) );
  OAI221XL U9518 ( .A0(n2221), .A1(n9487), .B0(n9551), .B1(n9374), .C0(n7225), 
        .Y(n2245) );
  OAI221XL U9519 ( .A0(n2221), .A1(n9484), .B0(n9542), .B1(n9374), .C0(n9623), 
        .Y(n2249) );
  NAND2X1 U9520 ( .A(n9710), .B(n9343), .Y(n145) );
  OAI21XL U9521 ( .A0(n9576), .A1(n2461), .B0(n7226), .Y(n2475) );
  OAI21XL U9522 ( .A0(n9567), .A1(n2461), .B0(n9636), .Y(n2479) );
  OAI21XL U9523 ( .A0(n351), .A1(n2461), .B0(n9632), .Y(n2483) );
  OAI21XL U9524 ( .A0(n9550), .A1(n2461), .B0(n7225), .Y(n2487) );
  OAI21XL U9525 ( .A0(n9540), .A1(n2461), .B0(n9623), .Y(n2492) );
  OAI21XL U9526 ( .A0(n7239), .A1(n1469), .B0(n7226), .Y(n1483) );
  OAI21XL U9527 ( .A0(n9567), .A1(n1469), .B0(n9638), .Y(n1487) );
  OAI21XL U9528 ( .A0(n9558), .A1(n1469), .B0(n9630), .Y(n1491) );
  OAI21XL U9529 ( .A0(n9551), .A1(n1469), .B0(n7225), .Y(n1495) );
  OAI21XL U9530 ( .A0(n9541), .A1(n1469), .B0(n9621), .Y(n1500) );
  OAI21XL U9531 ( .A0(n9578), .A1(n1782), .B0(n7226), .Y(n1796) );
  OAI21XL U9532 ( .A0(n9569), .A1(n1782), .B0(n9636), .Y(n1800) );
  OAI21XL U9533 ( .A0(n9558), .A1(n1782), .B0(n9630), .Y(n1804) );
  OAI21XL U9534 ( .A0(n9549), .A1(n1782), .B0(n7225), .Y(n1808) );
  OAI21XL U9535 ( .A0(n9541), .A1(n1782), .B0(n9621), .Y(n1813) );
  OAI21XL U9536 ( .A0(n9577), .A1(n1743), .B0(n7226), .Y(n1757) );
  OAI21XL U9537 ( .A0(n9567), .A1(n1743), .B0(n9638), .Y(n1761) );
  OAI21XL U9538 ( .A0(n9558), .A1(n1743), .B0(n9630), .Y(n1765) );
  OAI21XL U9539 ( .A0(n9550), .A1(n1743), .B0(n7225), .Y(n1769) );
  OAI21XL U9540 ( .A0(n9541), .A1(n1743), .B0(n9621), .Y(n1774) );
  OAI21XL U9541 ( .A0(n9576), .A1(n309), .B0(n7226), .Y(n334) );
  OAI21XL U9542 ( .A0(n9567), .A1(n309), .B0(n9636), .Y(n342) );
  OAI21XL U9543 ( .A0(n9558), .A1(n309), .B0(n9631), .Y(n350) );
  OAI21XL U9544 ( .A0(n9551), .A1(n309), .B0(n7225), .Y(n358) );
  OAI21XL U9545 ( .A0(n9540), .A1(n309), .B0(n9623), .Y(n371) );
  OAI21XL U9546 ( .A0(n9578), .A1(n382), .B0(n7226), .Y(n396) );
  OAI21XL U9547 ( .A0(n9569), .A1(n382), .B0(n9638), .Y(n400) );
  OAI21XL U9548 ( .A0(n9560), .A1(n382), .B0(n9632), .Y(n404) );
  OAI21XL U9549 ( .A0(n9550), .A1(n382), .B0(n7225), .Y(n408) );
  OAI21XL U9550 ( .A0(n9542), .A1(n382), .B0(n9623), .Y(n414) );
  OAI21XL U9551 ( .A0(n9578), .A1(n422), .B0(n7226), .Y(n436) );
  OAI21XL U9552 ( .A0(n9569), .A1(n422), .B0(n9638), .Y(n440) );
  OAI21XL U9553 ( .A0(n9560), .A1(n422), .B0(n9632), .Y(n444) );
  OAI21XL U9554 ( .A0(n9550), .A1(n422), .B0(n7225), .Y(n448) );
  OAI21XL U9555 ( .A0(n9542), .A1(n422), .B0(n9623), .Y(n454) );
  OAI21XL U9556 ( .A0(n9578), .A1(n462), .B0(n7226), .Y(n476) );
  OAI21XL U9557 ( .A0(n9569), .A1(n462), .B0(n9638), .Y(n480) );
  OAI21XL U9558 ( .A0(n9560), .A1(n462), .B0(n9632), .Y(n484) );
  OAI21XL U9559 ( .A0(n9550), .A1(n462), .B0(n7225), .Y(n488) );
  OAI21XL U9560 ( .A0(n9542), .A1(n462), .B0(n9623), .Y(n494) );
  OAI21XL U9561 ( .A0(n9578), .A1(n502), .B0(n7226), .Y(n516) );
  OAI21XL U9562 ( .A0(n9569), .A1(n502), .B0(n9638), .Y(n520) );
  OAI21XL U9563 ( .A0(n9560), .A1(n502), .B0(n9632), .Y(n524) );
  OAI21XL U9564 ( .A0(n9550), .A1(n502), .B0(n7225), .Y(n528) );
  OAI21XL U9565 ( .A0(n9542), .A1(n502), .B0(n9623), .Y(n534) );
  OAI21XL U9566 ( .A0(n9578), .A1(n542), .B0(n7226), .Y(n556) );
  OAI21XL U9567 ( .A0(n9569), .A1(n542), .B0(n9637), .Y(n560) );
  OAI21XL U9568 ( .A0(n9560), .A1(n542), .B0(n9631), .Y(n564) );
  OAI21XL U9569 ( .A0(n9550), .A1(n542), .B0(n7225), .Y(n568) );
  OAI21XL U9570 ( .A0(n9542), .A1(n542), .B0(n9622), .Y(n574) );
  OAI21XL U9571 ( .A0(n9578), .A1(n674), .B0(n7226), .Y(n688) );
  OAI21XL U9572 ( .A0(n9569), .A1(n674), .B0(n9638), .Y(n692) );
  OAI21XL U9573 ( .A0(n9560), .A1(n674), .B0(n9632), .Y(n696) );
  OAI21XL U9574 ( .A0(n9550), .A1(n674), .B0(n7225), .Y(n700) );
  OAI21XL U9575 ( .A0(n9542), .A1(n674), .B0(n9623), .Y(n707) );
  OAI21XL U9576 ( .A0(n9577), .A1(n715), .B0(n7226), .Y(n729) );
  OAI21XL U9577 ( .A0(n9568), .A1(n715), .B0(n9637), .Y(n733) );
  OAI21XL U9578 ( .A0(n9559), .A1(n715), .B0(n9631), .Y(n737) );
  OAI21XL U9579 ( .A0(n9549), .A1(n715), .B0(n7225), .Y(n741) );
  OAI21XL U9580 ( .A0(n9541), .A1(n715), .B0(n9622), .Y(n746) );
  OAI21XL U9581 ( .A0(n9578), .A1(n754), .B0(n7226), .Y(n768) );
  OAI21XL U9582 ( .A0(n9569), .A1(n754), .B0(n9638), .Y(n772) );
  OAI21XL U9583 ( .A0(n9560), .A1(n754), .B0(n9632), .Y(n776) );
  OAI21XL U9584 ( .A0(n9550), .A1(n754), .B0(n7225), .Y(n780) );
  OAI21XL U9585 ( .A0(n9542), .A1(n754), .B0(n9623), .Y(n785) );
  OAI21XL U9586 ( .A0(n9578), .A1(n793), .B0(n7226), .Y(n807) );
  OAI21XL U9587 ( .A0(n9569), .A1(n793), .B0(n9637), .Y(n811) );
  OAI21XL U9588 ( .A0(n9560), .A1(n793), .B0(n9631), .Y(n815) );
  OAI21XL U9589 ( .A0(n9550), .A1(n793), .B0(n7225), .Y(n819) );
  OAI21XL U9590 ( .A0(n9542), .A1(n793), .B0(n9622), .Y(n824) );
  OAI21XL U9591 ( .A0(n9577), .A1(n832), .B0(n7226), .Y(n846) );
  OAI21XL U9592 ( .A0(n9568), .A1(n832), .B0(n9638), .Y(n850) );
  OAI21XL U9593 ( .A0(n9559), .A1(n832), .B0(n9632), .Y(n854) );
  OAI21XL U9594 ( .A0(n9549), .A1(n832), .B0(n7225), .Y(n858) );
  OAI21XL U9595 ( .A0(n9540), .A1(n832), .B0(n9623), .Y(n863) );
  OAI21XL U9596 ( .A0(n9577), .A1(n871), .B0(n7226), .Y(n885) );
  OAI21XL U9597 ( .A0(n9568), .A1(n871), .B0(n9637), .Y(n889) );
  OAI21XL U9598 ( .A0(n9559), .A1(n871), .B0(n9630), .Y(n893) );
  OAI21XL U9599 ( .A0(n9549), .A1(n871), .B0(n7225), .Y(n897) );
  OAI21XL U9600 ( .A0(n9540), .A1(n871), .B0(n9621), .Y(n902) );
  OAI21XL U9601 ( .A0(n9577), .A1(n994), .B0(n7226), .Y(n1008) );
  OAI21XL U9602 ( .A0(n9568), .A1(n994), .B0(n9637), .Y(n1012) );
  OAI21XL U9603 ( .A0(n9559), .A1(n994), .B0(n9631), .Y(n1016) );
  OAI21XL U9604 ( .A0(n9549), .A1(n994), .B0(n7225), .Y(n1020) );
  OAI21XL U9605 ( .A0(n9541), .A1(n994), .B0(n9622), .Y(n1027) );
  OAI21XL U9606 ( .A0(n9577), .A1(n1035), .B0(n7226), .Y(n1049) );
  OAI21XL U9607 ( .A0(n9568), .A1(n1035), .B0(n9637), .Y(n1053) );
  OAI21XL U9608 ( .A0(n9559), .A1(n1035), .B0(n9631), .Y(n1057) );
  OAI21XL U9609 ( .A0(n9549), .A1(n1035), .B0(n7225), .Y(n1061) );
  OAI21XL U9610 ( .A0(n9540), .A1(n1035), .B0(n9622), .Y(n1066) );
  OAI21XL U9611 ( .A0(n9577), .A1(n1074), .B0(n7226), .Y(n1088) );
  OAI21XL U9612 ( .A0(n9568), .A1(n1074), .B0(n9637), .Y(n1092) );
  OAI21XL U9613 ( .A0(n9559), .A1(n1074), .B0(n9631), .Y(n1096) );
  OAI21XL U9614 ( .A0(n9549), .A1(n1074), .B0(n7225), .Y(n1100) );
  OAI21XL U9615 ( .A0(n9541), .A1(n1074), .B0(n9622), .Y(n1105) );
  OAI21XL U9616 ( .A0(n9577), .A1(n1113), .B0(n7226), .Y(n1127) );
  OAI21XL U9617 ( .A0(n9568), .A1(n1113), .B0(n9637), .Y(n1131) );
  OAI21XL U9618 ( .A0(n9559), .A1(n1113), .B0(n9631), .Y(n1135) );
  OAI21XL U9619 ( .A0(n9549), .A1(n1113), .B0(n7225), .Y(n1139) );
  OAI21XL U9620 ( .A0(n9541), .A1(n1113), .B0(n9622), .Y(n1144) );
  OAI21XL U9621 ( .A0(n9577), .A1(n1152), .B0(n7226), .Y(n1166) );
  OAI21XL U9622 ( .A0(n9568), .A1(n1152), .B0(n9637), .Y(n1170) );
  OAI21XL U9623 ( .A0(n9559), .A1(n1152), .B0(n9631), .Y(n1174) );
  OAI21XL U9624 ( .A0(n9549), .A1(n1152), .B0(n7225), .Y(n1178) );
  OAI21XL U9625 ( .A0(n9540), .A1(n1152), .B0(n9622), .Y(n1183) );
  OAI21XL U9626 ( .A0(n9577), .A1(n1191), .B0(n7226), .Y(n1205) );
  OAI21XL U9627 ( .A0(n9568), .A1(n1191), .B0(n9637), .Y(n1209) );
  OAI21XL U9628 ( .A0(n9559), .A1(n1191), .B0(n9631), .Y(n1213) );
  OAI21XL U9629 ( .A0(n9549), .A1(n1191), .B0(n7225), .Y(n1217) );
  OAI21XL U9630 ( .A0(n9541), .A1(n1191), .B0(n9622), .Y(n1222) );
  OAI21XL U9631 ( .A0(n9578), .A1(n1309), .B0(n7226), .Y(n1323) );
  OAI21XL U9632 ( .A0(n9568), .A1(n1309), .B0(n9637), .Y(n1327) );
  OAI21XL U9633 ( .A0(n9558), .A1(n1309), .B0(n9631), .Y(n1331) );
  OAI21XL U9634 ( .A0(n9549), .A1(n1309), .B0(n7225), .Y(n1335) );
  OAI21XL U9635 ( .A0(n9541), .A1(n1309), .B0(n9622), .Y(n1342) );
  OAI21XL U9636 ( .A0(n9578), .A1(n1350), .B0(n7226), .Y(n1364) );
  OAI21XL U9637 ( .A0(n9568), .A1(n1350), .B0(n9636), .Y(n1368) );
  OAI21XL U9638 ( .A0(n9558), .A1(n1350), .B0(n9630), .Y(n1372) );
  OAI21XL U9639 ( .A0(n9551), .A1(n1350), .B0(n7225), .Y(n1376) );
  OAI21XL U9640 ( .A0(n9541), .A1(n1350), .B0(n9621), .Y(n1381) );
  OAI21XL U9641 ( .A0(n9577), .A1(n1389), .B0(n7226), .Y(n1403) );
  OAI21XL U9642 ( .A0(n9568), .A1(n1389), .B0(n9637), .Y(n1407) );
  OAI21XL U9643 ( .A0(n9558), .A1(n1389), .B0(n9630), .Y(n1411) );
  OAI21XL U9644 ( .A0(n9549), .A1(n1389), .B0(n7225), .Y(n1415) );
  OAI21XL U9645 ( .A0(n9541), .A1(n1389), .B0(n9621), .Y(n1420) );
  OAI21XL U9646 ( .A0(n9577), .A1(n1508), .B0(n7226), .Y(n1522) );
  OAI21XL U9647 ( .A0(n9568), .A1(n1508), .B0(n9636), .Y(n1526) );
  OAI21XL U9648 ( .A0(n9558), .A1(n1508), .B0(n9630), .Y(n1530) );
  OAI21XL U9649 ( .A0(n9549), .A1(n1508), .B0(n7225), .Y(n1534) );
  OAI21XL U9650 ( .A0(n9541), .A1(n1508), .B0(n9621), .Y(n1539) );
  OAI21XL U9651 ( .A0(n9577), .A1(n1625), .B0(n7226), .Y(n1638) );
  OAI21XL U9652 ( .A0(n9568), .A1(n1625), .B0(n9637), .Y(n1642) );
  OAI21XL U9653 ( .A0(n9558), .A1(n1625), .B0(n9630), .Y(n1646) );
  OAI21XL U9654 ( .A0(n9549), .A1(n1625), .B0(n7225), .Y(n1650) );
  OAI21XL U9655 ( .A0(n9541), .A1(n1625), .B0(n9621), .Y(n1657) );
  OAI21XL U9656 ( .A0(n9578), .A1(n1665), .B0(n7226), .Y(n1679) );
  OAI21XL U9657 ( .A0(n9569), .A1(n1665), .B0(n9636), .Y(n1683) );
  OAI21XL U9658 ( .A0(n9558), .A1(n1665), .B0(n9630), .Y(n1687) );
  OAI21XL U9659 ( .A0(n9549), .A1(n1665), .B0(n7225), .Y(n1691) );
  OAI21XL U9660 ( .A0(n9541), .A1(n1665), .B0(n9621), .Y(n1696) );
  OAI21XL U9661 ( .A0(n9576), .A1(n1704), .B0(n7226), .Y(n1718) );
  OAI21XL U9662 ( .A0(n9568), .A1(n1704), .B0(n9637), .Y(n1722) );
  OAI21XL U9663 ( .A0(n9558), .A1(n1704), .B0(n9630), .Y(n1726) );
  OAI21XL U9664 ( .A0(n9549), .A1(n1704), .B0(n7225), .Y(n1730) );
  OAI21XL U9665 ( .A0(n9541), .A1(n1704), .B0(n9621), .Y(n1735) );
  OAI21XL U9666 ( .A0(n9576), .A1(n1823), .B0(n7226), .Y(n1837) );
  OAI21XL U9667 ( .A0(n9567), .A1(n1823), .B0(n9638), .Y(n1841) );
  OAI21XL U9668 ( .A0(n9558), .A1(n1823), .B0(n9630), .Y(n1845) );
  OAI21XL U9669 ( .A0(n9549), .A1(n1823), .B0(n7225), .Y(n1849) );
  OAI21XL U9670 ( .A0(n9541), .A1(n1823), .B0(n9621), .Y(n1854) );
  OAI21XL U9671 ( .A0(n9576), .A1(n1982), .B0(n7226), .Y(n1996) );
  OAI21XL U9672 ( .A0(n9567), .A1(n1982), .B0(n9636), .Y(n2000) );
  OAI21XL U9673 ( .A0(n9559), .A1(n1982), .B0(n9630), .Y(n2004) );
  OAI21XL U9674 ( .A0(n9550), .A1(n1982), .B0(n7225), .Y(n2008) );
  OAI21XL U9675 ( .A0(n9540), .A1(n1982), .B0(n9621), .Y(n2013) );
  OAI21XL U9676 ( .A0(n9577), .A1(n2021), .B0(n7226), .Y(n2035) );
  OAI21XL U9677 ( .A0(n9568), .A1(n2021), .B0(n9636), .Y(n2039) );
  OAI21XL U9678 ( .A0(n9559), .A1(n2021), .B0(n9631), .Y(n2043) );
  OAI21XL U9679 ( .A0(n9549), .A1(n2021), .B0(n7225), .Y(n2047) );
  OAI21XL U9680 ( .A0(n9541), .A1(n2021), .B0(n9622), .Y(n2052) );
  OAI21XL U9681 ( .A0(n9576), .A1(n2060), .B0(n7226), .Y(n2074) );
  OAI21XL U9682 ( .A0(n9567), .A1(n2060), .B0(n9636), .Y(n2078) );
  OAI21XL U9683 ( .A0(n9560), .A1(n2060), .B0(n9630), .Y(n2082) );
  OAI21XL U9684 ( .A0(n9549), .A1(n2060), .B0(n7225), .Y(n2086) );
  OAI21XL U9685 ( .A0(n9540), .A1(n2060), .B0(n9622), .Y(n2091) );
  OAI21XL U9686 ( .A0(n9576), .A1(n2099), .B0(n7226), .Y(n2113) );
  OAI21XL U9687 ( .A0(n9568), .A1(n2099), .B0(n9636), .Y(n2117) );
  OAI21XL U9688 ( .A0(n9560), .A1(n2099), .B0(n273), .Y(n2121) );
  OAI21XL U9689 ( .A0(n7238), .A1(n2099), .B0(n7225), .Y(n2125) );
  OAI21XL U9690 ( .A0(n9540), .A1(n2099), .B0(n287), .Y(n2134) );
  OAI21XL U9691 ( .A0(n9576), .A1(n2142), .B0(n7226), .Y(n2156) );
  OAI21XL U9692 ( .A0(n9567), .A1(n2142), .B0(n9636), .Y(n2160) );
  OAI21XL U9693 ( .A0(n9558), .A1(n2142), .B0(n9632), .Y(n2164) );
  OAI21XL U9694 ( .A0(n9551), .A1(n2142), .B0(n7225), .Y(n2168) );
  OAI21XL U9695 ( .A0(n9540), .A1(n2142), .B0(n9622), .Y(n2173) );
  OAI21XL U9696 ( .A0(n9576), .A1(n2260), .B0(n7226), .Y(n2273) );
  OAI21XL U9697 ( .A0(n9569), .A1(n2260), .B0(n9636), .Y(n2277) );
  OAI21XL U9698 ( .A0(n9558), .A1(n2260), .B0(n9632), .Y(n2281) );
  OAI21XL U9699 ( .A0(n7238), .A1(n2260), .B0(n7225), .Y(n2285) );
  OAI21XL U9700 ( .A0(n9540), .A1(n2260), .B0(n9621), .Y(n2293) );
  OAI21XL U9701 ( .A0(n9576), .A1(n2302), .B0(n7226), .Y(n2316) );
  OAI21XL U9702 ( .A0(n9568), .A1(n2302), .B0(n9636), .Y(n2320) );
  OAI21XL U9703 ( .A0(n351), .A1(n2302), .B0(n9630), .Y(n2324) );
  OAI21XL U9704 ( .A0(n9551), .A1(n2302), .B0(n7225), .Y(n2328) );
  OAI21XL U9705 ( .A0(n9540), .A1(n2302), .B0(n9623), .Y(n2333) );
  OAI21XL U9706 ( .A0(n9576), .A1(n2342), .B0(n7226), .Y(n2356) );
  OAI21XL U9707 ( .A0(n9567), .A1(n2342), .B0(n9636), .Y(n2360) );
  OAI21XL U9708 ( .A0(n351), .A1(n2342), .B0(n9631), .Y(n2364) );
  OAI21XL U9709 ( .A0(n9550), .A1(n2342), .B0(n7225), .Y(n2368) );
  OAI21XL U9710 ( .A0(n9540), .A1(n2342), .B0(n9621), .Y(n2373) );
  OAI21XL U9711 ( .A0(n9576), .A1(n2382), .B0(n7226), .Y(n2396) );
  OAI21XL U9712 ( .A0(n9567), .A1(n2382), .B0(n9636), .Y(n2400) );
  OAI21XL U9713 ( .A0(n351), .A1(n2382), .B0(n9631), .Y(n2404) );
  OAI21XL U9714 ( .A0(n9551), .A1(n2382), .B0(n7225), .Y(n2408) );
  OAI21XL U9715 ( .A0(n9540), .A1(n2382), .B0(n9621), .Y(n2414) );
  OAI21XL U9716 ( .A0(n9570), .A1(n9347), .B0(n7226), .Y(n2516) );
  OAI21XL U9717 ( .A0(n9562), .A1(n9347), .B0(n9637), .Y(n2520) );
  OAI21XL U9718 ( .A0(n9552), .A1(n9347), .B0(n9631), .Y(n2524) );
  OAI21XL U9719 ( .A0(n9543), .A1(n9347), .B0(n7225), .Y(n2528) );
  OAI21XL U9720 ( .A0(n9534), .A1(n9347), .B0(n9622), .Y(n2533) );
  BUFX4 U9721 ( .A(n8940), .Y(n8942) );
  CLKBUFX3 U9722 ( .A(n8939), .Y(n8943) );
  CLKBUFX3 U9723 ( .A(n8939), .Y(n8944) );
  BUFX4 U9724 ( .A(n8956), .Y(n8958) );
  BUFX4 U9725 ( .A(n8955), .Y(n8959) );
  CLKBUFX3 U9726 ( .A(n8964), .Y(n8960) );
  CLKBUFX3 U9727 ( .A(n8955), .Y(n8961) );
  CLKBUFX3 U9728 ( .A(n8964), .Y(n8963) );
  CLKBUFX3 U9729 ( .A(n266), .Y(n9636) );
  CLKBUFX3 U9730 ( .A(n9144), .Y(n9147) );
  CLKBUFX3 U9731 ( .A(n9145), .Y(n9148) );
  CLKBUFX3 U9732 ( .A(n9145), .Y(n9146) );
  CLKBUFX3 U9733 ( .A(n110), .Y(n9444) );
  OAI21XL U9734 ( .A0(n9665), .A1(n7226), .B0(n9640), .Y(n110) );
  CLKBUFX3 U9735 ( .A(n113), .Y(n9442) );
  OAI21XL U9736 ( .A0(n9665), .A1(n9636), .B0(n9633), .Y(n113) );
  CLKBUFX3 U9737 ( .A(n116), .Y(n9440) );
  OAI21XL U9738 ( .A0(n9666), .A1(n9630), .B0(n9627), .Y(n116) );
  CLKBUFX3 U9739 ( .A(n8956), .Y(n8957) );
  CLKBUFX3 U9740 ( .A(n8940), .Y(n8941) );
  CLKBUFX3 U9741 ( .A(n8932), .Y(n8934) );
  CLKBUFX3 U9742 ( .A(n8931), .Y(n8938) );
  CLKBUFX3 U9743 ( .A(n8932), .Y(n8935) );
  CLKINVX1 U9744 ( .A(n9512), .Y(n8925) );
  CLKINVX1 U9745 ( .A(n9516), .Y(n9125) );
  OAI221XL U9746 ( .A0(n1428), .A1(n9505), .B0(n9604), .B1(n1429), .C0(n9659), 
        .Y(n1424) );
  OAI221XL U9747 ( .A0(n1428), .A1(n9502), .B0(n9596), .B1(n1429), .C0(n9653), 
        .Y(n1432) );
  OAI221XL U9748 ( .A0(n1428), .A1(n9499), .B0(n9587), .B1(n1429), .C0(n9647), 
        .Y(n1436) );
  OAI221XL U9749 ( .A0(n1941), .A1(n9505), .B0(n9604), .B1(n1942), .C0(n9659), 
        .Y(n1937) );
  OAI221XL U9750 ( .A0(n1941), .A1(n9502), .B0(n9596), .B1(n1942), .C0(n9653), 
        .Y(n1945) );
  OAI221XL U9751 ( .A0(n1941), .A1(n9499), .B0(n9587), .B1(n1942), .C0(n9647), 
        .Y(n1949) );
  OAI221XL U9752 ( .A0(n2422), .A1(n9505), .B0(n9605), .B1(n2423), .C0(n235), 
        .Y(n2418) );
  OAI221XL U9753 ( .A0(n2422), .A1(n9502), .B0(n9594), .B1(n2423), .C0(n9652), 
        .Y(n2426) );
  OAI221XL U9754 ( .A0(n2422), .A1(n9499), .B0(n9586), .B1(n2423), .C0(n9646), 
        .Y(n2430) );
  OAI221XL U9755 ( .A0(n2422), .A1(n9498), .B0(n9576), .B1(n2423), .C0(n7226), 
        .Y(n2434) );
  OAI221XL U9756 ( .A0(n1902), .A1(n9505), .B0(n9605), .B1(n1903), .C0(n9657), 
        .Y(n1898) );
  OAI221XL U9757 ( .A0(n1902), .A1(n9502), .B0(n9596), .B1(n1903), .C0(n9652), 
        .Y(n1906) );
  OAI221XL U9758 ( .A0(n1902), .A1(n9499), .B0(n9586), .B1(n1903), .C0(n9646), 
        .Y(n1910) );
  OAI221XL U9759 ( .A0(n1902), .A1(n9497), .B0(n9577), .B1(n1903), .C0(n7226), 
        .Y(n1914) );
  OAI221XL U9760 ( .A0(n626), .A1(n9505), .B0(n9605), .B1(n9422), .C0(n9659), 
        .Y(n621) );
  OAI221XL U9761 ( .A0(n626), .A1(n9502), .B0(n8417), .B1(n9422), .C0(n9653), 
        .Y(n630) );
  OAI221XL U9762 ( .A0(n626), .A1(n9499), .B0(n9585), .B1(n9422), .C0(n9647), 
        .Y(n635) );
  OAI221XL U9763 ( .A0(n950), .A1(n9505), .B0(n9604), .B1(n9412), .C0(n9659), 
        .Y(n946) );
  OAI221XL U9764 ( .A0(n950), .A1(n9502), .B0(n9596), .B1(n9412), .C0(n9653), 
        .Y(n954) );
  OAI221XL U9765 ( .A0(n950), .A1(n9499), .B0(n9587), .B1(n9412), .C0(n9647), 
        .Y(n958) );
  OAI221XL U9766 ( .A0(n1270), .A1(n9505), .B0(n9604), .B1(n9402), .C0(n9659), 
        .Y(n1266) );
  OAI221XL U9767 ( .A0(n1270), .A1(n9502), .B0(n9596), .B1(n9402), .C0(n9653), 
        .Y(n1274) );
  OAI221XL U9768 ( .A0(n1270), .A1(n9499), .B0(n9587), .B1(n9402), .C0(n9647), 
        .Y(n1278) );
  OAI221XL U9769 ( .A0(n1587), .A1(n9505), .B0(n9604), .B1(n9392), .C0(n9659), 
        .Y(n1583) );
  OAI221XL U9770 ( .A0(n1587), .A1(n9502), .B0(n9596), .B1(n9392), .C0(n9653), 
        .Y(n1591) );
  OAI221XL U9771 ( .A0(n1587), .A1(n9499), .B0(n9587), .B1(n9392), .C0(n9647), 
        .Y(n1595) );
  OAI221XL U9772 ( .A0(n2221), .A1(n9505), .B0(n9605), .B1(n9374), .C0(n9659), 
        .Y(n2217) );
  OAI221XL U9773 ( .A0(n2221), .A1(n9502), .B0(n9594), .B1(n9374), .C0(n9653), 
        .Y(n2225) );
  OAI221XL U9774 ( .A0(n2221), .A1(n9499), .B0(n9586), .B1(n9374), .C0(n9647), 
        .Y(n2229) );
  OAI21XL U9775 ( .A0(n9603), .A1(n2461), .B0(n9657), .Y(n2460) );
  OAI21XL U9776 ( .A0(n9594), .A1(n2461), .B0(n9651), .Y(n2467) );
  OAI21XL U9777 ( .A0(n9587), .A1(n2461), .B0(n9645), .Y(n2471) );
  OAI21XL U9778 ( .A0(n9604), .A1(n1469), .B0(n9658), .Y(n1468) );
  OAI21XL U9779 ( .A0(n9594), .A1(n1469), .B0(n9652), .Y(n1475) );
  OAI21XL U9780 ( .A0(n9585), .A1(n1469), .B0(n9646), .Y(n1479) );
  OAI21XL U9781 ( .A0(n308), .A1(n1782), .B0(n9658), .Y(n1781) );
  OAI21XL U9782 ( .A0(n9594), .A1(n1782), .B0(n9652), .Y(n1788) );
  OAI21XL U9783 ( .A0(n9585), .A1(n1782), .B0(n9646), .Y(n1792) );
  OAI21XL U9784 ( .A0(n308), .A1(n1743), .B0(n9658), .Y(n1742) );
  OAI21XL U9785 ( .A0(n9594), .A1(n1743), .B0(n9652), .Y(n1749) );
  OAI21XL U9786 ( .A0(n9585), .A1(n1743), .B0(n9646), .Y(n1753) );
  OAI21XL U9787 ( .A0(n9603), .A1(n309), .B0(n9657), .Y(n307) );
  OAI21XL U9788 ( .A0(n9595), .A1(n309), .B0(n9651), .Y(n318) );
  OAI21XL U9789 ( .A0(n9585), .A1(n309), .B0(n9645), .Y(n326) );
  OAI21XL U9790 ( .A0(n9604), .A1(n382), .B0(n9659), .Y(n381) );
  OAI21XL U9791 ( .A0(n9596), .A1(n382), .B0(n9653), .Y(n388) );
  OAI21XL U9792 ( .A0(n9587), .A1(n382), .B0(n9647), .Y(n392) );
  OAI21XL U9793 ( .A0(n9604), .A1(n422), .B0(n9659), .Y(n421) );
  OAI21XL U9794 ( .A0(n9596), .A1(n422), .B0(n9653), .Y(n428) );
  OAI21XL U9795 ( .A0(n9587), .A1(n422), .B0(n9647), .Y(n432) );
  OAI21XL U9796 ( .A0(n9604), .A1(n462), .B0(n9659), .Y(n461) );
  OAI21XL U9797 ( .A0(n9596), .A1(n462), .B0(n9653), .Y(n468) );
  OAI21XL U9798 ( .A0(n9587), .A1(n462), .B0(n9647), .Y(n472) );
  OAI21XL U9799 ( .A0(n9604), .A1(n502), .B0(n9659), .Y(n501) );
  OAI21XL U9800 ( .A0(n9596), .A1(n502), .B0(n9653), .Y(n508) );
  OAI21XL U9801 ( .A0(n9587), .A1(n502), .B0(n9647), .Y(n512) );
  OAI21XL U9802 ( .A0(n9604), .A1(n542), .B0(n9658), .Y(n541) );
  OAI21XL U9803 ( .A0(n9596), .A1(n542), .B0(n9653), .Y(n548) );
  OAI21XL U9804 ( .A0(n9587), .A1(n542), .B0(n9647), .Y(n552) );
  OAI21XL U9805 ( .A0(n9604), .A1(n674), .B0(n9659), .Y(n673) );
  OAI21XL U9806 ( .A0(n9596), .A1(n674), .B0(n9653), .Y(n680) );
  OAI21XL U9807 ( .A0(n9587), .A1(n674), .B0(n9647), .Y(n684) );
  OAI21XL U9808 ( .A0(n9605), .A1(n715), .B0(n235), .Y(n714) );
  OAI21XL U9809 ( .A0(n9595), .A1(n715), .B0(n245), .Y(n721) );
  OAI21XL U9810 ( .A0(n9586), .A1(n715), .B0(n9646), .Y(n725) );
  OAI21XL U9811 ( .A0(n9604), .A1(n754), .B0(n9659), .Y(n753) );
  OAI21XL U9812 ( .A0(n9596), .A1(n754), .B0(n9653), .Y(n760) );
  OAI21XL U9813 ( .A0(n9587), .A1(n754), .B0(n9647), .Y(n764) );
  OAI21XL U9814 ( .A0(n9604), .A1(n793), .B0(n9658), .Y(n792) );
  OAI21XL U9815 ( .A0(n9596), .A1(n793), .B0(n9652), .Y(n799) );
  OAI21XL U9816 ( .A0(n9587), .A1(n793), .B0(n252), .Y(n803) );
  OAI21XL U9817 ( .A0(n9605), .A1(n832), .B0(n9659), .Y(n831) );
  OAI21XL U9818 ( .A0(n9595), .A1(n832), .B0(n9653), .Y(n838) );
  OAI21XL U9819 ( .A0(n9586), .A1(n832), .B0(n9647), .Y(n842) );
  OAI21XL U9820 ( .A0(n9605), .A1(n871), .B0(n9658), .Y(n870) );
  OAI21XL U9821 ( .A0(n9595), .A1(n871), .B0(n9652), .Y(n877) );
  OAI21XL U9822 ( .A0(n9586), .A1(n871), .B0(n9646), .Y(n881) );
  OAI21XL U9823 ( .A0(n9605), .A1(n994), .B0(n9658), .Y(n993) );
  OAI21XL U9824 ( .A0(n9595), .A1(n994), .B0(n245), .Y(n1000) );
  OAI21XL U9825 ( .A0(n9586), .A1(n994), .B0(n9645), .Y(n1004) );
  OAI21XL U9826 ( .A0(n9605), .A1(n1035), .B0(n9658), .Y(n1034) );
  OAI21XL U9827 ( .A0(n9595), .A1(n1035), .B0(n9652), .Y(n1041) );
  OAI21XL U9828 ( .A0(n9586), .A1(n1035), .B0(n9646), .Y(n1045) );
  OAI21XL U9829 ( .A0(n9605), .A1(n1074), .B0(n9658), .Y(n1073) );
  OAI21XL U9830 ( .A0(n9595), .A1(n1074), .B0(n245), .Y(n1080) );
  OAI21XL U9831 ( .A0(n9586), .A1(n1074), .B0(n252), .Y(n1084) );
  OAI21XL U9832 ( .A0(n9605), .A1(n1113), .B0(n9658), .Y(n1112) );
  OAI21XL U9833 ( .A0(n9595), .A1(n1113), .B0(n9651), .Y(n1119) );
  OAI21XL U9834 ( .A0(n9586), .A1(n1113), .B0(n9646), .Y(n1123) );
  OAI21XL U9835 ( .A0(n9605), .A1(n1152), .B0(n235), .Y(n1151) );
  OAI21XL U9836 ( .A0(n9595), .A1(n1152), .B0(n9652), .Y(n1158) );
  OAI21XL U9837 ( .A0(n9586), .A1(n1152), .B0(n9646), .Y(n1162) );
  OAI21XL U9838 ( .A0(n9603), .A1(n1191), .B0(n235), .Y(n1190) );
  OAI21XL U9839 ( .A0(n9595), .A1(n1191), .B0(n245), .Y(n1197) );
  OAI21XL U9840 ( .A0(n9586), .A1(n1191), .B0(n9646), .Y(n1201) );
  OAI21XL U9841 ( .A0(n9604), .A1(n1309), .B0(n235), .Y(n1308) );
  OAI21XL U9842 ( .A0(n9595), .A1(n1309), .B0(n9652), .Y(n1315) );
  OAI21XL U9843 ( .A0(n9585), .A1(n1309), .B0(n252), .Y(n1319) );
  OAI21XL U9844 ( .A0(n308), .A1(n1350), .B0(n9658), .Y(n1349) );
  OAI21XL U9845 ( .A0(n9594), .A1(n1350), .B0(n9652), .Y(n1356) );
  OAI21XL U9846 ( .A0(n9585), .A1(n1350), .B0(n9646), .Y(n1360) );
  OAI21XL U9847 ( .A0(n308), .A1(n1389), .B0(n9658), .Y(n1388) );
  OAI21XL U9848 ( .A0(n9595), .A1(n1389), .B0(n9652), .Y(n1395) );
  OAI21XL U9849 ( .A0(n9585), .A1(n1389), .B0(n9646), .Y(n1399) );
  OAI21XL U9850 ( .A0(n9604), .A1(n1508), .B0(n9658), .Y(n1507) );
  OAI21XL U9851 ( .A0(n9594), .A1(n1508), .B0(n9652), .Y(n1514) );
  OAI21XL U9852 ( .A0(n9585), .A1(n1508), .B0(n9646), .Y(n1518) );
  OAI21XL U9853 ( .A0(n9604), .A1(n1625), .B0(n9658), .Y(n1624) );
  OAI21XL U9854 ( .A0(n9596), .A1(n1625), .B0(n9652), .Y(n1630) );
  OAI21XL U9855 ( .A0(n9585), .A1(n1625), .B0(n9646), .Y(n1634) );
  OAI21XL U9856 ( .A0(n9605), .A1(n1665), .B0(n9658), .Y(n1664) );
  OAI21XL U9857 ( .A0(n9594), .A1(n1665), .B0(n9652), .Y(n1671) );
  OAI21XL U9858 ( .A0(n9585), .A1(n1665), .B0(n9646), .Y(n1675) );
  OAI21XL U9859 ( .A0(n9604), .A1(n1704), .B0(n9658), .Y(n1703) );
  OAI21XL U9860 ( .A0(n9595), .A1(n1704), .B0(n9652), .Y(n1710) );
  OAI21XL U9861 ( .A0(n9585), .A1(n1704), .B0(n9646), .Y(n1714) );
  OAI21XL U9862 ( .A0(n9605), .A1(n1823), .B0(n9658), .Y(n1822) );
  OAI21XL U9863 ( .A0(n9595), .A1(n1823), .B0(n9652), .Y(n1829) );
  OAI21XL U9864 ( .A0(n9585), .A1(n1823), .B0(n9646), .Y(n1833) );
  OAI21XL U9865 ( .A0(n9603), .A1(n1982), .B0(n9657), .Y(n1981) );
  OAI21XL U9866 ( .A0(n8417), .A1(n1982), .B0(n9651), .Y(n1988) );
  OAI21XL U9867 ( .A0(n9586), .A1(n1982), .B0(n9645), .Y(n1992) );
  OAI21XL U9868 ( .A0(n308), .A1(n2021), .B0(n9657), .Y(n2020) );
  OAI21XL U9869 ( .A0(n9595), .A1(n2021), .B0(n9651), .Y(n2027) );
  OAI21XL U9870 ( .A0(n9586), .A1(n2021), .B0(n252), .Y(n2031) );
  OAI21XL U9871 ( .A0(n9603), .A1(n2060), .B0(n9657), .Y(n2059) );
  OAI21XL U9872 ( .A0(n8417), .A1(n2060), .B0(n9651), .Y(n2066) );
  OAI21XL U9873 ( .A0(n9587), .A1(n2060), .B0(n9645), .Y(n2070) );
  OAI21XL U9874 ( .A0(n9603), .A1(n2099), .B0(n9657), .Y(n2098) );
  OAI21XL U9875 ( .A0(n9595), .A1(n2099), .B0(n9651), .Y(n2105) );
  OAI21XL U9876 ( .A0(n9587), .A1(n2099), .B0(n9645), .Y(n2109) );
  OAI21XL U9877 ( .A0(n9603), .A1(n2142), .B0(n9657), .Y(n2141) );
  OAI21XL U9878 ( .A0(n9594), .A1(n2142), .B0(n9651), .Y(n2148) );
  OAI21XL U9879 ( .A0(n9585), .A1(n2142), .B0(n9645), .Y(n2152) );
  OAI21XL U9880 ( .A0(n9603), .A1(n2260), .B0(n9657), .Y(n2259) );
  OAI21XL U9881 ( .A0(n9595), .A1(n2260), .B0(n9651), .Y(n2265) );
  OAI21XL U9882 ( .A0(n9587), .A1(n2260), .B0(n9645), .Y(n2269) );
  OAI21XL U9883 ( .A0(n9603), .A1(n2302), .B0(n9657), .Y(n2301) );
  OAI21XL U9884 ( .A0(n9596), .A1(n2302), .B0(n9651), .Y(n2308) );
  OAI21XL U9885 ( .A0(n9585), .A1(n2302), .B0(n9645), .Y(n2312) );
  OAI21XL U9886 ( .A0(n9603), .A1(n2342), .B0(n9657), .Y(n2341) );
  OAI21XL U9887 ( .A0(n9594), .A1(n2342), .B0(n9651), .Y(n2348) );
  OAI21XL U9888 ( .A0(n9587), .A1(n2342), .B0(n9645), .Y(n2352) );
  OAI21XL U9889 ( .A0(n9603), .A1(n2382), .B0(n9657), .Y(n2381) );
  OAI21XL U9890 ( .A0(n8417), .A1(n2382), .B0(n9651), .Y(n2388) );
  OAI21XL U9891 ( .A0(n9586), .A1(n2382), .B0(n9645), .Y(n2392) );
  OAI21XL U9892 ( .A0(n9597), .A1(n9347), .B0(n9658), .Y(n2500) );
  OAI21XL U9893 ( .A0(n9588), .A1(n9347), .B0(n245), .Y(n2508) );
  OAI21XL U9894 ( .A0(n9579), .A1(n9347), .B0(n9645), .Y(n2512) );
  CLKBUFX3 U9895 ( .A(n9138), .Y(n9139) );
  CLKBUFX3 U9896 ( .A(n9138), .Y(n8929) );
  CLKBUFX3 U9897 ( .A(n9152), .Y(n8962) );
  CLKBUFX3 U9898 ( .A(n9127), .Y(n8919) );
  CLKBUFX3 U9899 ( .A(n235), .Y(n9657) );
  CLKBUFX3 U9900 ( .A(n245), .Y(n9651) );
  CLKBUFX3 U9901 ( .A(n9145), .Y(n9149) );
  CLKBUFX3 U9902 ( .A(n9144), .Y(n9150) );
  CLKBUFX3 U9903 ( .A(n9143), .Y(n9151) );
  CLKBUFX3 U9904 ( .A(n9511), .Y(n8928) );
  CLKBUFX3 U9905 ( .A(n100), .Y(n9450) );
  OAI21XL U9906 ( .A0(n9665), .A1(n9657), .B0(n9654), .Y(n100) );
  CLKBUFX3 U9907 ( .A(n104), .Y(n9448) );
  OAI21XL U9908 ( .A0(n9665), .A1(n9651), .B0(n9649), .Y(n104) );
  CLKBUFX3 U9909 ( .A(n107), .Y(n9446) );
  OAI21XL U9910 ( .A0(n9665), .A1(n9645), .B0(n9643), .Y(n107) );
  CLKBUFX3 U9911 ( .A(n8931), .Y(n8937) );
  CLKINVX1 U9912 ( .A(n9512), .Y(n8924) );
  CLKINVX1 U9913 ( .A(n9356), .Y(n9733) );
  CLKINVX1 U9914 ( .A(n9355), .Y(n9732) );
  CLKINVX1 U9915 ( .A(n9354), .Y(n9731) );
  CLKINVX1 U9916 ( .A(n9353), .Y(n9730) );
  CLKINVX1 U9917 ( .A(n9352), .Y(n9729) );
  CLKINVX1 U9918 ( .A(n9351), .Y(n9728) );
  CLKINVX1 U9919 ( .A(n9350), .Y(n9727) );
  CLKINVX1 U9920 ( .A(n9346), .Y(n9726) );
  CLKBUFX3 U9921 ( .A(n320), .Y(n9591) );
  CLKBUFX3 U9922 ( .A(n328), .Y(n9582) );
  CLKBUFX3 U9923 ( .A(n336), .Y(n9573) );
  CLKBUFX3 U9924 ( .A(n344), .Y(n9564) );
  CLKBUFX3 U9925 ( .A(n345), .Y(n9561) );
  CLKBUFX3 U9926 ( .A(n8417), .Y(n9594) );
  CLKBUFX3 U9927 ( .A(n308), .Y(n9605) );
  CLKBUFX3 U9928 ( .A(n7237), .Y(n9567) );
  CLKBUFX3 U9929 ( .A(n7238), .Y(n9551) );
  CLKINVX1 U9930 ( .A(n9435), .Y(n9718) );
  CLKINVX1 U9931 ( .A(n9449), .Y(n9725) );
  CLKINVX1 U9932 ( .A(n9447), .Y(n9724) );
  CLKINVX1 U9933 ( .A(n9445), .Y(n9723) );
  CLKINVX1 U9934 ( .A(n9443), .Y(n9722) );
  CLKINVX1 U9935 ( .A(n9441), .Y(n9721) );
  CLKINVX1 U9936 ( .A(n9439), .Y(n9720) );
  CLKINVX1 U9937 ( .A(n9437), .Y(n9719) );
  AOI2BB2X2 U9938 ( .B0(n9610), .B1(n9789), .A0N(n9616), .A1N(n9414), .Y(n583)
         );
  AOI2BB2X2 U9939 ( .B0(n9609), .B1(n9757), .A0N(n9615), .A1N(n9781), .Y(n1470) );
  NOR2BX2 U9940 ( .AN(n9433), .B(n9421), .Y(n233) );
  OA22X2 U9941 ( .A0(n9616), .A1(n9347), .B0(n9611), .B1(n7236), .Y(n2504) );
  OA22X2 U9942 ( .A0(n9616), .A1(n9521), .B0(n9612), .B1(n9523), .Y(n1902) );
  OA22X2 U9943 ( .A0(n9616), .A1(n2183), .B0(n9612), .B1(n9521), .Y(n2182) );
  OA22X2 U9944 ( .A0(n9616), .A1(n9404), .B0(n9611), .B1(n9533), .Y(n911) );
  OA22X2 U9945 ( .A0(n9616), .A1(n9394), .B0(n9611), .B1(n9531), .Y(n1231) );
  OA22X2 U9946 ( .A0(n9616), .A1(n9384), .B0(n9611), .B1(n9527), .Y(n1548) );
  OA22X2 U9947 ( .A0(n9616), .A1(n9376), .B0(n9611), .B1(n9525), .Y(n1863) );
  NAND3X2 U9948 ( .A(n7236), .B(n9345), .C(n9347), .Y(n2503) );
  NAND3X2 U9949 ( .A(n9524), .B(n9522), .C(n9520), .Y(n1903) );
  INVX3 U9950 ( .A(n9424), .Y(n9790) );
  CLKBUFX3 U9951 ( .A(n625), .Y(n9532) );
  CLKBUFX3 U9952 ( .A(n949), .Y(n9530) );
  CLKBUFX3 U9953 ( .A(n1269), .Y(n9526) );
  CLKBUFX3 U9954 ( .A(n1586), .Y(n9524) );
  CLKBUFX3 U9955 ( .A(n1901), .Y(n9520) );
  INVX3 U9956 ( .A(n9617), .Y(n9614) );
  INVX3 U9957 ( .A(n9414), .Y(n9749) );
  CLKBUFX3 U9958 ( .A(n9812), .Y(n9505) );
  CLKBUFX3 U9959 ( .A(n9811), .Y(n9502) );
  CLKBUFX3 U9960 ( .A(n9810), .Y(n9499) );
  CLKBUFX3 U9961 ( .A(n9807), .Y(n9490) );
  CLKBUFX3 U9962 ( .A(n9806), .Y(n9487) );
  CLKBUFX3 U9963 ( .A(n9805), .Y(n9484) );
  CLKBUFX3 U9964 ( .A(n9812), .Y(n9507) );
  CLKBUFX3 U9965 ( .A(n9812), .Y(n9506) );
  CLKBUFX3 U9966 ( .A(n9811), .Y(n9504) );
  CLKBUFX3 U9967 ( .A(n9810), .Y(n9501) );
  CLKBUFX3 U9968 ( .A(n9809), .Y(n9498) );
  CLKBUFX3 U9969 ( .A(n9808), .Y(n9495) );
  CLKBUFX3 U9970 ( .A(n9807), .Y(n9492) );
  CLKBUFX3 U9971 ( .A(n9806), .Y(n9489) );
  CLKBUFX3 U9972 ( .A(n9805), .Y(n9486) );
  CLKBUFX3 U9973 ( .A(n9811), .Y(n9503) );
  CLKBUFX3 U9974 ( .A(n9810), .Y(n9500) );
  CLKBUFX3 U9975 ( .A(n9809), .Y(n9497) );
  CLKBUFX3 U9976 ( .A(n9808), .Y(n9494) );
  CLKBUFX3 U9977 ( .A(n9806), .Y(n9488) );
  CLKBUFX3 U9978 ( .A(n9805), .Y(n9485) );
  CLKBUFX3 U9979 ( .A(n9809), .Y(n9496) );
  CLKBUFX3 U9980 ( .A(n9808), .Y(n9493) );
  CLKBUFX3 U9981 ( .A(n9807), .Y(n9491) );
  CLKINVX1 U9982 ( .A(n9421), .Y(n9789) );
  CLKBUFX3 U9983 ( .A(n625), .Y(n9533) );
  CLKBUFX3 U9984 ( .A(n949), .Y(n9531) );
  CLKBUFX3 U9985 ( .A(n1269), .Y(n9527) );
  CLKBUFX3 U9986 ( .A(n1586), .Y(n9525) );
  CLKBUFX3 U9987 ( .A(n1901), .Y(n9521) );
  AOI2BB2X2 U9988 ( .B0(n9610), .B1(n9776), .A0N(n9615), .A1N(n9529), .Y(n1114) );
  AOI2BB2X2 U9989 ( .B0(n9609), .B1(n9787), .A0N(n9614), .A1N(n9523), .Y(n1626) );
  AOI2BB2X2 U9990 ( .B0(n9608), .B1(n9763), .A0N(n9614), .A1N(n9519), .Y(n2100) );
  NAND2X2 U9991 ( .A(n9434), .B(n9796), .Y(n241) );
  INVX3 U9992 ( .A(n2183), .Y(n9768) );
  INVX3 U9993 ( .A(n9404), .Y(n9774) );
  INVX3 U9994 ( .A(n9394), .Y(n9756) );
  INVX3 U9995 ( .A(n9384), .Y(n9783) );
  INVX3 U9996 ( .A(n9376), .Y(n9762) );
  INVX3 U9997 ( .A(n9612), .Y(n9607) );
  CLKBUFX3 U9998 ( .A(n218), .Y(n9434) );
  NOR2X1 U9999 ( .A(n9614), .B(n9664), .Y(n218) );
  INVX3 U10000 ( .A(n9611), .Y(n9608) );
  INVX3 U10001 ( .A(n9611), .Y(n9609) );
  CLKBUFX3 U10002 ( .A(n219), .Y(n9433) );
  NOR2X1 U10003 ( .A(n9611), .B(n9664), .Y(n219) );
  INVX3 U10004 ( .A(n9611), .Y(n9610) );
  INVX3 U10005 ( .A(n9613), .Y(n9616) );
  INVX3 U10006 ( .A(n9665), .Y(n9663) );
  INVX3 U10007 ( .A(n9665), .Y(n9662) );
  INVX3 U10008 ( .A(n9665), .Y(n9661) );
  CLKBUFX3 U10009 ( .A(n9332), .Y(n9325) );
  CLKBUFX3 U10010 ( .A(n9332), .Y(n9327) );
  CLKBUFX3 U10011 ( .A(n9332), .Y(n9326) );
  CLKBUFX3 U10012 ( .A(n9332), .Y(n9328) );
  CLKBUFX3 U10013 ( .A(n9332), .Y(n9329) );
  CLKBUFX3 U10014 ( .A(n9332), .Y(n9331) );
  CLKBUFX3 U10015 ( .A(n9332), .Y(n9330) );
  CLKBUFX3 U10016 ( .A(N1656), .Y(n9316) );
  CLKBUFX3 U10017 ( .A(N1656), .Y(n9315) );
  CLKBUFX3 U10018 ( .A(N1656), .Y(n9314) );
  NOR2X2 U10019 ( .A(n9665), .B(n9423), .Y(n623) );
  NOR2X2 U10020 ( .A(n9665), .B(n9403), .Y(n1268) );
  NOR2X2 U10021 ( .A(n9666), .B(n9393), .Y(n1585) );
  NOR2X2 U10022 ( .A(n9665), .B(n9383), .Y(n1900) );
  NOR2X2 U10023 ( .A(n9665), .B(n9375), .Y(n2219) );
  NAND2X2 U10024 ( .A(n9663), .B(n703), .Y(n669) );
  NAND2X2 U10025 ( .A(n9663), .B(n744), .Y(n710) );
  NAND2X2 U10026 ( .A(n9663), .B(n783), .Y(n749) );
  NAND2X2 U10027 ( .A(n9662), .B(n822), .Y(n788) );
  NAND2X2 U10028 ( .A(n9662), .B(n861), .Y(n827) );
  NAND2X2 U10029 ( .A(n9662), .B(n900), .Y(n866) );
  NAND2X2 U10030 ( .A(n9662), .B(n939), .Y(n905) );
  NAND2X2 U10031 ( .A(n9662), .B(n1023), .Y(n989) );
  NAND2X2 U10032 ( .A(n9662), .B(n1064), .Y(n1030) );
  NAND2X2 U10033 ( .A(n9662), .B(n1103), .Y(n1069) );
  NAND2X2 U10034 ( .A(n9662), .B(n1142), .Y(n1108) );
  NAND2X2 U10035 ( .A(n9662), .B(n1181), .Y(n1147) );
  NAND2X2 U10036 ( .A(n9662), .B(n1220), .Y(n1186) );
  NAND2X2 U10037 ( .A(n9662), .B(n1259), .Y(n1225) );
  NAND2X2 U10038 ( .A(n9661), .B(n1653), .Y(n1620) );
  NAND2X2 U10039 ( .A(n9662), .B(n1694), .Y(n1660) );
  NAND2X2 U10040 ( .A(n9661), .B(n1733), .Y(n1699) );
  NAND2X2 U10041 ( .A(n9662), .B(n1772), .Y(n1738) );
  NAND2X2 U10042 ( .A(n9661), .B(n1811), .Y(n1777) );
  NAND2X2 U10043 ( .A(n9661), .B(n1852), .Y(n1818) );
  NAND2X2 U10044 ( .A(n9661), .B(n1891), .Y(n1857) );
  NAND2X2 U10045 ( .A(n9662), .B(n1338), .Y(n1304) );
  NAND2X2 U10046 ( .A(n9661), .B(n1379), .Y(n1345) );
  NAND2X2 U10047 ( .A(n9663), .B(n1418), .Y(n1384) );
  NAND2X2 U10048 ( .A(n9662), .B(n1498), .Y(n1464) );
  NAND2X2 U10049 ( .A(n9663), .B(n1537), .Y(n1503) );
  NAND2X2 U10050 ( .A(n9663), .B(n1576), .Y(n1542) );
  NAND2X2 U10051 ( .A(n9661), .B(n2050), .Y(n2016) );
  NAND2X2 U10052 ( .A(n9661), .B(n2089), .Y(n2055) );
  NAND2X2 U10053 ( .A(n9661), .B(n2128), .Y(n2094) );
  NAND2X2 U10054 ( .A(n9661), .B(n2171), .Y(n2137) );
  NAND2X2 U10055 ( .A(n9661), .B(n2210), .Y(n2176) );
  NAND2X2 U10056 ( .A(n9661), .B(n2288), .Y(n2255) );
  NAND2X2 U10057 ( .A(n9661), .B(n2371), .Y(n2336) );
  NAND2X2 U10058 ( .A(n9661), .B(n2411), .Y(n2376) );
  NAND2X2 U10059 ( .A(n9661), .B(n2490), .Y(n2456) );
  NAND2X2 U10060 ( .A(n9661), .B(n2531), .Y(n2495) );
  NAND2X2 U10061 ( .A(n9663), .B(n364), .Y(n302) );
  NAND2X2 U10062 ( .A(n9663), .B(n411), .Y(n377) );
  NAND2X2 U10063 ( .A(n9663), .B(n451), .Y(n417) );
  NAND2X2 U10064 ( .A(n9663), .B(n491), .Y(n457) );
  NAND2X2 U10065 ( .A(n9663), .B(n611), .Y(n577) );
  INVX3 U10066 ( .A(n9458), .Y(n9668) );
  INVX3 U10067 ( .A(n703), .Y(n9708) );
  INVX3 U10068 ( .A(n744), .Y(n9702) );
  INVX3 U10069 ( .A(n783), .Y(n9695) );
  INVX3 U10070 ( .A(n822), .Y(n9688) );
  INVX3 U10071 ( .A(n861), .Y(n9715) );
  INVX3 U10072 ( .A(n900), .Y(n9682) );
  INVX3 U10073 ( .A(n939), .Y(n9675) );
  INVX3 U10074 ( .A(n1023), .Y(n9707) );
  INVX3 U10075 ( .A(n1064), .Y(n9701) );
  INVX3 U10076 ( .A(n1103), .Y(n9694) );
  INVX3 U10077 ( .A(n1142), .Y(n9687) );
  INVX3 U10078 ( .A(n1181), .Y(n9714) );
  INVX3 U10079 ( .A(n1220), .Y(n9681) );
  INVX3 U10080 ( .A(n1259), .Y(n9674) );
  INVX3 U10081 ( .A(n1653), .Y(n9705) );
  INVX3 U10082 ( .A(n1694), .Y(n9699) );
  INVX3 U10083 ( .A(n1733), .Y(n9692) );
  INVX3 U10084 ( .A(n1772), .Y(n9686) );
  INVX3 U10085 ( .A(n1811), .Y(n9712) );
  INVX3 U10086 ( .A(n1852), .Y(n9679) );
  INVX3 U10087 ( .A(n1891), .Y(n9672) );
  INVX3 U10088 ( .A(n1338), .Y(n9706) );
  INVX3 U10089 ( .A(n1379), .Y(n9700) );
  INVX3 U10090 ( .A(n1418), .Y(n9693) );
  INVX3 U10091 ( .A(n1498), .Y(n9713) );
  INVX3 U10092 ( .A(n1537), .Y(n9680) );
  INVX3 U10093 ( .A(n1576), .Y(n9673) );
  INVX3 U10094 ( .A(n2011), .Y(n9698) );
  INVX3 U10095 ( .A(n2050), .Y(n9691) );
  INVX3 U10096 ( .A(n2089), .Y(n9685) );
  INVX3 U10097 ( .A(n2128), .Y(n9711) );
  INVX3 U10098 ( .A(n2171), .Y(n9678) );
  INVX3 U10099 ( .A(n2210), .Y(n9671) );
  INVX3 U10100 ( .A(n2288), .Y(n9704) );
  INVX3 U10101 ( .A(n2331), .Y(n9697) );
  INVX3 U10102 ( .A(n2371), .Y(n9690) );
  INVX3 U10103 ( .A(n2411), .Y(n9684) );
  INVX3 U10104 ( .A(n2490), .Y(n9677) );
  INVX3 U10105 ( .A(n2531), .Y(n9670) );
  INVX3 U10106 ( .A(n364), .Y(n9709) );
  INVX3 U10107 ( .A(n411), .Y(n9703) );
  INVX3 U10108 ( .A(n451), .Y(n9696) );
  INVX3 U10109 ( .A(n491), .Y(n9689) );
  INVX3 U10110 ( .A(n531), .Y(n9716) );
  INVX3 U10111 ( .A(n571), .Y(n9683) );
  INVX3 U10112 ( .A(n611), .Y(n9676) );
  CLKINVX1 U10113 ( .A(n230), .Y(n9710) );
  CLKBUFX3 U10114 ( .A(n188), .Y(n9453) );
  OA22X1 U10115 ( .A0(n159), .A1(n199), .B0(n200), .B1(n145), .Y(n188) );
  CLKBUFX3 U10116 ( .A(n9153), .Y(n9145) );
  CLKBUFX3 U10117 ( .A(n8930), .Y(n8939) );
  CLKBUFX3 U10118 ( .A(n9153), .Y(n8956) );
  CLKBUFX3 U10119 ( .A(n8930), .Y(n8940) );
  CLKBUFX3 U10120 ( .A(n8964), .Y(n8955) );
  CLKBUFX3 U10121 ( .A(n8954), .Y(n8931) );
  CLKBUFX3 U10122 ( .A(n8954), .Y(n8932) );
  NOR2X2 U10123 ( .A(n9413), .B(n9664), .Y(n948) );
  NOR2X2 U10124 ( .A(n9382), .B(n9665), .Y(n1939) );
  CLKBUFX3 U10125 ( .A(n236), .Y(n9654) );
  CLKBUFX3 U10126 ( .A(n9648), .Y(n9649) );
  CLKBUFX3 U10127 ( .A(n9642), .Y(n9643) );
  CLKBUFX3 U10128 ( .A(n9639), .Y(n9640) );
  CLKBUFX3 U10129 ( .A(n267), .Y(n9633) );
  CLKBUFX3 U10130 ( .A(n274), .Y(n9627) );
  CLKBUFX3 U10131 ( .A(n281), .Y(n9625) );
  CLKBUFX3 U10132 ( .A(n288), .Y(n9618) );
  CLKBUFX3 U10133 ( .A(n9655), .Y(n9656) );
  CLKBUFX3 U10134 ( .A(n9649), .Y(n9650) );
  CLKBUFX3 U10135 ( .A(n9643), .Y(n9644) );
  CLKBUFX3 U10136 ( .A(n9640), .Y(n9641) );
  CLKBUFX3 U10137 ( .A(n274), .Y(n9629) );
  CLKBUFX3 U10138 ( .A(n9624), .Y(n9626) );
  CLKBUFX3 U10139 ( .A(n9618), .Y(n9620) );
  CLKBUFX3 U10140 ( .A(n236), .Y(n9655) );
  CLKBUFX3 U10141 ( .A(n267), .Y(n9634) );
  CLKBUFX3 U10142 ( .A(n274), .Y(n9628) );
  CLKBUFX3 U10143 ( .A(n288), .Y(n9619) );
  CLKBUFX3 U10144 ( .A(n8922), .Y(n9136) );
  CLKBUFX3 U10145 ( .A(n9634), .Y(n9635) );
  CLKBUFX3 U10146 ( .A(n252), .Y(n9645) );
  CLKBUFX3 U10147 ( .A(n9153), .Y(n9144) );
  CLKBUFX3 U10148 ( .A(n9152), .Y(n9143) );
  AO22X1 U10149 ( .A0(n9434), .A1(N7387), .B0(n9433), .B1(n8436), .Y(n128) );
  AO22X1 U10150 ( .A0(n9434), .A1(N7386), .B0(n9433), .B1(n8437), .Y(n131) );
  AO22X1 U10151 ( .A0(n9434), .A1(N7385), .B0(n9433), .B1(n8434), .Y(n133) );
  AO22X1 U10152 ( .A0(n9434), .A1(N7384), .B0(n9433), .B1(n8435), .Y(n135) );
  AO22X1 U10153 ( .A0(n9434), .A1(N7383), .B0(n9433), .B1(n8442), .Y(n137) );
  AO22X1 U10154 ( .A0(n9434), .A1(N7382), .B0(n9433), .B1(n8443), .Y(n139) );
  AO22X1 U10155 ( .A0(n9434), .A1(N7381), .B0(n9433), .B1(n8444), .Y(n141) );
  AO22X1 U10156 ( .A0(n9434), .A1(N7380), .B0(n9433), .B1(n8445), .Y(n143) );
  NAND2X1 U10157 ( .A(n8436), .B(n9613), .Y(n310) );
  NAND2X1 U10158 ( .A(n8437), .B(n9613), .Y(n320) );
  NAND2X1 U10159 ( .A(n8434), .B(n9613), .Y(n328) );
  NAND2X1 U10160 ( .A(n8435), .B(n9613), .Y(n336) );
  NAND2X1 U10161 ( .A(n8442), .B(n9617), .Y(n344) );
  NAND2X1 U10162 ( .A(n8443), .B(n9613), .Y(n352) );
  NAND2X1 U10163 ( .A(n8444), .B(n9617), .Y(n360) );
  NAND2X1 U10164 ( .A(n8445), .B(n9613), .Y(n373) );
  AO22X1 U10165 ( .A0(n292), .A1(N7388), .B0(n9608), .B1(n8419), .Y(n8432) );
  CLKINVX1 U10166 ( .A(n8432), .Y(n308) );
  NAND2X1 U10167 ( .A(n8437), .B(n9610), .Y(n321) );
  NAND2X1 U10168 ( .A(n8434), .B(n9610), .Y(n329) );
  NAND2X1 U10169 ( .A(n8435), .B(n9610), .Y(n337) );
  NAND2X1 U10170 ( .A(n8442), .B(n9610), .Y(n345) );
  NAND2X1 U10171 ( .A(n8443), .B(n9610), .Y(n353) );
  NAND2X1 U10172 ( .A(n8444), .B(n9610), .Y(n361) );
  NAND2X1 U10173 ( .A(n8445), .B(n9609), .Y(n374) );
  NAND2X1 U10174 ( .A(n8436), .B(n9610), .Y(n313) );
  CLKBUFX3 U10175 ( .A(n101), .Y(n9449) );
  CLKBUFX3 U10176 ( .A(n105), .Y(n9447) );
  AO22X1 U10177 ( .A0(n9433), .A1(n8420), .B0(n9434), .B1(n8418), .Y(n105) );
  CLKBUFX3 U10178 ( .A(n108), .Y(n9445) );
  AO22X1 U10179 ( .A0(n9433), .A1(n7227), .B0(n9434), .B1(n7233), .Y(n108) );
  CLKBUFX3 U10180 ( .A(n111), .Y(n9443) );
  AO22X1 U10181 ( .A0(n9433), .A1(n7234), .B0(n9434), .B1(N7391), .Y(n111) );
  CLKBUFX3 U10182 ( .A(n114), .Y(n9441) );
  AO22X1 U10183 ( .A0(n9433), .A1(n7228), .B0(n9434), .B1(N7392), .Y(n114) );
  CLKBUFX3 U10184 ( .A(n117), .Y(n9439) );
  AO22X1 U10185 ( .A0(n9433), .A1(n7229), .B0(n9434), .B1(N7393), .Y(n117) );
  CLKBUFX3 U10186 ( .A(n120), .Y(n9437) );
  AO22X1 U10187 ( .A0(n9433), .A1(n7230), .B0(n9434), .B1(n7235), .Y(n120) );
  CLKBUFX3 U10188 ( .A(n123), .Y(n9435) );
  AO22X1 U10189 ( .A0(n9433), .A1(n7231), .B0(n9434), .B1(N7395), .Y(n123) );
  CLKBUFX3 U10190 ( .A(n632), .Y(n9355) );
  AOI22X1 U10191 ( .A0(n8418), .A1(n9607), .B0(n8420), .B1(n9613), .Y(n632) );
  CLKBUFX3 U10192 ( .A(n637), .Y(n9354) );
  AOI22X1 U10193 ( .A0(n7233), .A1(n9607), .B0(n7227), .B1(n9617), .Y(n637) );
  CLKBUFX3 U10194 ( .A(n642), .Y(n9353) );
  AOI22X1 U10195 ( .A0(N7391), .A1(n9607), .B0(n7234), .B1(n9613), .Y(n642) );
  CLKBUFX3 U10196 ( .A(n647), .Y(n9352) );
  AOI22X1 U10197 ( .A0(N7392), .A1(n9607), .B0(n7228), .B1(n9613), .Y(n647) );
  CLKBUFX3 U10198 ( .A(n652), .Y(n9351) );
  AOI22X1 U10199 ( .A0(N7393), .A1(n9607), .B0(n7229), .B1(n9613), .Y(n652) );
  CLKBUFX3 U10200 ( .A(n657), .Y(n9350) );
  AOI22X1 U10201 ( .A0(n7235), .A1(n9607), .B0(n7230), .B1(n9617), .Y(n657) );
  CLKBUFX3 U10202 ( .A(n662), .Y(n9346) );
  AOI22X1 U10203 ( .A0(N7395), .A1(n9607), .B0(n7231), .B1(n9613), .Y(n662) );
  CLKBUFX3 U10204 ( .A(n624), .Y(n9356) );
  INVX3 U10205 ( .A(n9512), .Y(n9137) );
  AO22X1 U10206 ( .A0(n9613), .A1(N7393), .B0(n9608), .B1(n7229), .Y(n8433) );
  CLKINVX1 U10207 ( .A(n8433), .Y(n351) );
  CLKBUFX3 U10208 ( .A(n9152), .Y(n9142) );
  OAI21X2 U10209 ( .A0(n2211), .A1(n9373), .B0(n9349), .Y(n1973) );
  OAI21X2 U10210 ( .A0(n9344), .A1(n9391), .B0(n9349), .Y(n1340) );
  OAI21X2 U10211 ( .A0(n2294), .A1(n2211), .B0(n9349), .Y(n2290) );
  AOI2BB2X2 U10212 ( .B0(n9610), .B1(n9790), .A0N(n9615), .A1N(n9415), .Y(n543) );
  AOI2BB2X2 U10213 ( .B0(n9607), .B1(n9749), .A0N(n9615), .A1N(n9405), .Y(n872) );
  NAND2X1 U10214 ( .A(n667), .B(n9411), .Y(n625) );
  NAND2X1 U10215 ( .A(n9401), .B(n667), .Y(n949) );
  NAND2X1 U10216 ( .A(n9391), .B(n667), .Y(n1269) );
  NAND2X1 U10217 ( .A(n9344), .B(n667), .Y(n1586) );
  NAND2X1 U10218 ( .A(n9373), .B(n667), .Y(n1901) );
  INVX3 U10219 ( .A(n9430), .Y(n9796) );
  NOR2X1 U10220 ( .A(n667), .B(n617), .Y(n228) );
  BUFX4 U10221 ( .A(n584), .Y(n9414) );
  NAND2X1 U10222 ( .A(n9411), .B(n617), .Y(n584) );
  CLKBUFX3 U10223 ( .A(n229), .Y(n9343) );
  NOR3X1 U10224 ( .A(n9512), .B(n9514), .C(n9510), .Y(n229) );
  BUFX4 U10225 ( .A(n296), .Y(n9421) );
  NAND2X1 U10226 ( .A(n667), .B(n9343), .Y(n296) );
  NAND2X1 U10227 ( .A(n617), .B(n9343), .Y(n217) );
  CLKBUFX3 U10228 ( .A(n9613), .Y(n9617) );
  CLKBUFX3 U10229 ( .A(n9660), .Y(n9666) );
  CLKBUFX3 U10230 ( .A(n1775), .Y(n9386) );
  NOR2X1 U10231 ( .A(n9782), .B(n9813), .Y(n1775) );
  CLKBUFX3 U10232 ( .A(n627), .Y(n9422) );
  NAND3X1 U10233 ( .A(n9421), .B(n9420), .C(n9532), .Y(n627) );
  CLKBUFX3 U10234 ( .A(n1271), .Y(n9402) );
  NAND3X1 U10235 ( .A(n9530), .B(n9400), .C(n9526), .Y(n1271) );
  CLKBUFX3 U10236 ( .A(n240), .Y(n9431) );
  NAND2X1 U10237 ( .A(n9421), .B(n9430), .Y(n240) );
  CLKBUFX3 U10238 ( .A(n1588), .Y(n9392) );
  NAND3X1 U10239 ( .A(n9526), .B(n9390), .C(n9524), .Y(n1588) );
  CLKBUFX3 U10240 ( .A(n2222), .Y(n9374) );
  NAND3X1 U10241 ( .A(n9520), .B(n9371), .C(n7236), .Y(n2222) );
  CLKBUFX3 U10242 ( .A(n951), .Y(n9412) );
  NAND3X1 U10243 ( .A(n9532), .B(n9410), .C(n9530), .Y(n951) );
  OAI21X2 U10244 ( .A0(n9343), .A1(n9411), .B0(n9349), .Y(n367) );
  OAI21X2 U10245 ( .A0(n9401), .A1(n9411), .B0(n9349), .Y(n705) );
  OAI21X2 U10246 ( .A0(n9391), .A1(n9401), .B0(n9349), .Y(n1025) );
  OAI21X2 U10247 ( .A0(n9344), .A1(n9373), .B0(n9349), .Y(n1655) );
  AOI2BB2X2 U10248 ( .B0(n9610), .B1(n9795), .A0N(n9614), .A1N(n9420), .Y(n311) );
  AOI2BB2X2 U10249 ( .B0(n9610), .B1(n9794), .A0N(n9616), .A1N(n9419), .Y(n383) );
  AOI2BB2X2 U10250 ( .B0(n9610), .B1(n9793), .A0N(n9616), .A1N(n9418), .Y(n423) );
  AOI2BB2X2 U10251 ( .B0(n9610), .B1(n9792), .A0N(n9616), .A1N(n9417), .Y(n463) );
  AOI2BB2X2 U10252 ( .B0(n9610), .B1(n9791), .A0N(n9616), .A1N(n9416), .Y(n503) );
  AOI2BB2X2 U10253 ( .B0(n9607), .B1(n9754), .A0N(n9615), .A1N(n9410), .Y(n675) );
  AOI2BB2X2 U10254 ( .B0(n293), .B1(n9753), .A0N(n9615), .A1N(n9409), .Y(n716)
         );
  AOI2BB2X2 U10255 ( .B0(n9607), .B1(n9752), .A0N(n9615), .A1N(n9408), .Y(n755) );
  AOI2BB2X2 U10256 ( .B0(n9607), .B1(n9751), .A0N(n9615), .A1N(n9407), .Y(n794) );
  AOI2BB2X2 U10257 ( .B0(n9607), .B1(n9750), .A0N(n9615), .A1N(n9406), .Y(n833) );
  AOI2BB2X2 U10258 ( .B0(n9609), .B1(n9779), .A0N(n9615), .A1N(n9400), .Y(n995) );
  AOI2BB2X2 U10259 ( .B0(n9606), .B1(n9778), .A0N(n9615), .A1N(n9399), .Y(
        n1036) );
  AOI2BB2X2 U10260 ( .B0(n9606), .B1(n9777), .A0N(n9615), .A1N(n9398), .Y(
        n1075) );
  AOI2BB2X2 U10261 ( .B0(n293), .B1(n9775), .A0N(n9615), .A1N(n9396), .Y(n1153) );
  AOI2BB2X2 U10262 ( .B0(n9609), .B1(n9774), .A0N(n9615), .A1N(n9395), .Y(
        n1192) );
  AOI2BB2X2 U10263 ( .B0(n9609), .B1(n9760), .A0N(n9615), .A1N(n9390), .Y(
        n1310) );
  AOI2BB2X2 U10264 ( .B0(n9609), .B1(n9759), .A0N(n9615), .A1N(n9389), .Y(
        n1351) );
  AOI2BB2X2 U10265 ( .B0(n9609), .B1(n9756), .A0N(n9614), .A1N(n9385), .Y(
        n1509) );
  AOI2BB2X2 U10266 ( .B0(n9609), .B1(n9786), .A0N(n9614), .A1N(n9381), .Y(
        n1666) );
  AOI2BB2X2 U10267 ( .B0(n9609), .B1(n9785), .A0N(n9614), .A1N(n9380), .Y(
        n1705) );
  AOI2BB2X2 U10268 ( .B0(n9609), .B1(n9386), .A0N(n9614), .A1N(n9379), .Y(
        n1744) );
  AOI2BB2X2 U10269 ( .B0(n9608), .B1(n9784), .A0N(n9614), .A1N(n9378), .Y(
        n1783) );
  AOI2BB2X2 U10270 ( .B0(n9608), .B1(n9783), .A0N(n9614), .A1N(n9377), .Y(
        n1824) );
  AOI2BB2X2 U10271 ( .B0(n9608), .B1(n9766), .A0N(n9614), .A1N(n9369), .Y(
        n1983) );
  AOI2BB2X2 U10272 ( .B0(n9608), .B1(n9765), .A0N(n9614), .A1N(n9366), .Y(
        n2022) );
  AOI2BB2X2 U10273 ( .B0(n9608), .B1(n9764), .A0N(n9614), .A1N(n9363), .Y(
        n2061) );
  AOI2BB2X2 U10274 ( .B0(n9608), .B1(n9762), .A0N(n9614), .A1N(n9358), .Y(
        n2143) );
  OA22X2 U10275 ( .A0(n9611), .A1(n9345), .B0(n9616), .B1(n9359), .Y(n2463) );
  OA22X2 U10276 ( .A0(n9616), .A1(n9388), .B0(n9611), .B1(n9529), .Y(n1390) );
  OA22X2 U10277 ( .A0(n9612), .A1(n9369), .B0(n9616), .B1(n9372), .Y(n2261) );
  OA22X2 U10278 ( .A0(n9611), .A1(n9366), .B0(n9616), .B1(n9370), .Y(n2304) );
  OA22X2 U10279 ( .A0(n9611), .A1(n9363), .B0(n9616), .B1(n9367), .Y(n2344) );
  OA22X2 U10280 ( .A0(n9611), .A1(n9519), .B0(n9616), .B1(n9364), .Y(n2384) );
  NAND2X2 U10281 ( .A(n2211), .B(n617), .Y(n2183) );
  NAND3X2 U10282 ( .A(n9396), .B(n9528), .C(n9387), .Y(n1429) );
  NAND3X2 U10283 ( .A(n9381), .B(n9522), .C(n9371), .Y(n1942) );
  NAND3X2 U10284 ( .A(n9358), .B(n9518), .C(n9361), .Y(n2423) );
  AND2X2 U10285 ( .A(n2535), .B(n9510), .Y(n2294) );
  NAND2X2 U10286 ( .A(n2211), .B(n617), .Y(n9345) );
  INVX3 U10287 ( .A(n9369), .Y(n9772) );
  INVX3 U10288 ( .A(n9366), .Y(n9771) );
  INVX3 U10289 ( .A(n9363), .Y(n9770) );
  INVX3 U10290 ( .A(n9429), .Y(n9795) );
  INVX3 U10291 ( .A(n9428), .Y(n9794) );
  INVX3 U10292 ( .A(n9427), .Y(n9793) );
  INVX3 U10293 ( .A(n9426), .Y(n9792) );
  INVX3 U10294 ( .A(n9425), .Y(n9791) );
  BUFX4 U10295 ( .A(n912), .Y(n9404) );
  NAND2X1 U10296 ( .A(n9401), .B(n617), .Y(n912) );
  BUFX4 U10297 ( .A(n1232), .Y(n9394) );
  NAND2X1 U10298 ( .A(n9391), .B(n617), .Y(n1232) );
  BUFX4 U10299 ( .A(n1549), .Y(n9384) );
  NAND2X1 U10300 ( .A(n9344), .B(n617), .Y(n1549) );
  BUFX4 U10301 ( .A(n1864), .Y(n9376) );
  NAND2X1 U10302 ( .A(n9373), .B(n617), .Y(n1864) );
  CLKBUFX3 U10303 ( .A(n7247), .Y(n9528) );
  CLKBUFX3 U10304 ( .A(n7248), .Y(n9518) );
  INVX3 U10305 ( .A(n9410), .Y(n9780) );
  INVX3 U10306 ( .A(n9390), .Y(n9788) );
  INVX3 U10307 ( .A(n9371), .Y(n9773) );
  INVX3 U10308 ( .A(n9420), .Y(n9755) );
  INVX3 U10309 ( .A(n9400), .Y(n9761) );
  CLKINVX1 U10310 ( .A(n9344), .Y(n9782) );
  INVX3 U10311 ( .A(n9358), .Y(n9769) );
  INVX3 U10312 ( .A(n9419), .Y(n9754) );
  INVX3 U10313 ( .A(n9418), .Y(n9753) );
  INVX3 U10314 ( .A(n9417), .Y(n9752) );
  INVX3 U10315 ( .A(n9416), .Y(n9751) );
  INVX3 U10316 ( .A(n9415), .Y(n9750) );
  INVX3 U10317 ( .A(n9409), .Y(n9779) );
  INVX3 U10318 ( .A(n9408), .Y(n9778) );
  INVX3 U10319 ( .A(n9407), .Y(n9777) );
  INVX3 U10320 ( .A(n9406), .Y(n9776) );
  INVX3 U10321 ( .A(n9405), .Y(n9775) );
  INVX3 U10322 ( .A(n9399), .Y(n9760) );
  INVX3 U10323 ( .A(n9398), .Y(n9759) );
  INVX3 U10324 ( .A(n9396), .Y(n9758) );
  INVX3 U10325 ( .A(n9395), .Y(n9757) );
  INVX3 U10326 ( .A(n9389), .Y(n9787) );
  INVX3 U10327 ( .A(n9387), .Y(n9785) );
  INVX3 U10328 ( .A(n9385), .Y(n9784) );
  INVX3 U10329 ( .A(n9381), .Y(n9767) );
  INVX3 U10330 ( .A(n9380), .Y(n9766) );
  INVX3 U10331 ( .A(n9379), .Y(n9765) );
  INVX3 U10332 ( .A(n9378), .Y(n9764) );
  INVX3 U10333 ( .A(n9377), .Y(n9763) );
  INVX3 U10334 ( .A(n9388), .Y(n9786) );
  CLKBUFX3 U10335 ( .A(n9612), .Y(n9611) );
  CLKBUFX3 U10336 ( .A(n2501), .Y(n9347) );
  NAND2X1 U10337 ( .A(n2294), .B(n617), .Y(n2501) );
  CLKBUFX3 U10338 ( .A(n7248), .Y(n9519) );
  CLKBUFX3 U10339 ( .A(n7245), .Y(n9523) );
  CLKBUFX3 U10340 ( .A(n7247), .Y(n9529) );
  CLKBUFX3 U10341 ( .A(n9660), .Y(n9665) );
  NAND2X1 U10342 ( .A(n2569), .B(n9459), .Y(n2570) );
  CLKBUFX3 U10343 ( .A(n9669), .Y(n9459) );
  CLKBUFX3 U10344 ( .A(N1659), .Y(n9335) );
  CLKBUFX3 U10345 ( .A(N1659), .Y(n9336) );
  CLKBUFX3 U10346 ( .A(n9334), .Y(n9333) );
  NAND2BX2 U10347 ( .AN(n161), .B(n2129), .Y(n412) );
  NAND2BX2 U10348 ( .AN(n174), .B(n2129), .Y(n452) );
  NAND2BX2 U10349 ( .AN(n213), .B(n2129), .Y(n572) );
  NAND2BX2 U10350 ( .AN(n228), .B(n2129), .Y(n612) );
  MX4X1 U10351 ( .A(n8984), .B(n8974), .C(n8979), .D(n8969), .S0(n9136), .S1(
        n9137), .Y(N7387) );
  MX4X1 U10352 ( .A(n8973), .B(n8971), .C(n8972), .D(n8970), .S0(n9139), .S1(
        n9140), .Y(n8974) );
  MX4X1 U10353 ( .A(n8968), .B(n8966), .C(n8967), .D(n8965), .S0(n9139), .S1(
        n9140), .Y(n8969) );
  MX4X1 U10354 ( .A(n8983), .B(n8981), .C(n8982), .D(n8980), .S0(n9139), .S1(
        n9140), .Y(n8984) );
  CLKBUFX3 U10355 ( .A(n98), .Y(n9458) );
  AOI32X1 U10356 ( .A0(N1677), .A1(n9669), .A2(n96), .B0(n9710), .B1(n9796), 
        .Y(n98) );
  NAND2BX1 U10357 ( .AN(n200), .B(n2129), .Y(n532) );
  NAND2BX1 U10358 ( .AN(n144), .B(n2129), .Y(n368) );
  NAND2BX1 U10359 ( .AN(n187), .B(n2129), .Y(n492) );
  OAI22X1 U10360 ( .A0(n8106), .A1(n365), .B0(n367), .B1(n412), .Y(n411) );
  OAI22X1 U10361 ( .A0(n8263), .A1(n365), .B0(n367), .B1(n452), .Y(n451) );
  OAI22X1 U10362 ( .A0(n8329), .A1(n365), .B0(n367), .B1(n612), .Y(n611) );
  OAI22X1 U10363 ( .A0(n8106), .A1(n704), .B0(n412), .B1(n705), .Y(n744) );
  OAI22X1 U10364 ( .A0(n8263), .A1(n704), .B0(n452), .B1(n705), .Y(n783) );
  OAI22X1 U10365 ( .A0(n8312), .A1(n704), .B0(n572), .B1(n705), .Y(n900) );
  OAI22X1 U10366 ( .A0(n8329), .A1(n704), .B0(n612), .B1(n705), .Y(n939) );
  OAI22X1 U10367 ( .A0(n8106), .A1(n7807), .B0(n412), .B1(n1025), .Y(n1064) );
  OAI22X1 U10368 ( .A0(n8263), .A1(n7807), .B0(n452), .B1(n1025), .Y(n1103) );
  OAI22X1 U10369 ( .A0(n8312), .A1(n7807), .B0(n572), .B1(n1025), .Y(n1220) );
  OAI22X1 U10370 ( .A0(n8329), .A1(n7807), .B0(n612), .B1(n1025), .Y(n1259) );
  OAI22X1 U10371 ( .A0(n8106), .A1(n1339), .B0(n412), .B1(n1340), .Y(n1379) );
  OAI22X1 U10372 ( .A0(n8263), .A1(n1339), .B0(n452), .B1(n1340), .Y(n1418) );
  OAI22X1 U10373 ( .A0(n8312), .A1(n1339), .B0(n572), .B1(n1340), .Y(n1537) );
  OAI22X1 U10374 ( .A0(n8329), .A1(n1339), .B0(n612), .B1(n1340), .Y(n1576) );
  OAI22X1 U10375 ( .A0(n8106), .A1(n8187), .B0(n412), .B1(n1655), .Y(n1694) );
  OAI22X1 U10376 ( .A0(n8263), .A1(n8187), .B0(n452), .B1(n1655), .Y(n1733) );
  OAI22X1 U10377 ( .A0(n8312), .A1(n8187), .B0(n572), .B1(n1655), .Y(n1852) );
  OAI22X1 U10378 ( .A0(n8329), .A1(n8187), .B0(n612), .B1(n1655), .Y(n1891) );
  OAI22X1 U10379 ( .A0(n160), .A1(n1974), .B0(n412), .B1(n1973), .Y(n2011) );
  OAI22X1 U10380 ( .A0(n8263), .A1(n1974), .B0(n452), .B1(n1973), .Y(n2050) );
  OAI22X1 U10381 ( .A0(n8312), .A1(n1974), .B0(n572), .B1(n1973), .Y(n2171) );
  OAI22X1 U10382 ( .A0(n8329), .A1(n1974), .B0(n612), .B1(n1973), .Y(n2210) );
  OAI22X1 U10383 ( .A0(n9340), .A1(n8263), .B0(n452), .B1(n2290), .Y(n2371) );
  OAI22X1 U10384 ( .A0(n9340), .A1(n8312), .B0(n572), .B1(n2290), .Y(n2490) );
  OAI22X1 U10385 ( .A0(n9340), .A1(n8329), .B0(n612), .B1(n2290), .Y(n2531) );
  OAI22X1 U10386 ( .A0(n366), .A1(n704), .B0(n368), .B1(n705), .Y(n703) );
  OAI22X1 U10387 ( .A0(n186), .A1(n704), .B0(n492), .B1(n705), .Y(n822) );
  OAI22X1 U10388 ( .A0(n199), .A1(n704), .B0(n532), .B1(n705), .Y(n861) );
  OAI22X1 U10389 ( .A0(n366), .A1(n7807), .B0(n368), .B1(n1025), .Y(n1023) );
  OAI22X1 U10390 ( .A0(n186), .A1(n7807), .B0(n492), .B1(n1025), .Y(n1142) );
  OAI22X1 U10391 ( .A0(n199), .A1(n7807), .B0(n532), .B1(n1025), .Y(n1181) );
  OAI22X1 U10392 ( .A0(n366), .A1(n8187), .B0(n368), .B1(n1655), .Y(n1653) );
  OAI22X1 U10393 ( .A0(n186), .A1(n8187), .B0(n492), .B1(n1655), .Y(n1772) );
  OAI22X1 U10394 ( .A0(n199), .A1(n8187), .B0(n532), .B1(n1655), .Y(n1811) );
  OAI22X1 U10395 ( .A0(n365), .A1(n366), .B0(n367), .B1(n368), .Y(n364) );
  OAI22X1 U10396 ( .A0(n186), .A1(n365), .B0(n367), .B1(n492), .Y(n491) );
  OAI22X1 U10397 ( .A0(n366), .A1(n1339), .B0(n368), .B1(n1340), .Y(n1338) );
  OAI22X1 U10398 ( .A0(n199), .A1(n1339), .B0(n532), .B1(n1340), .Y(n1498) );
  OAI22X1 U10399 ( .A0(n186), .A1(n1974), .B0(n492), .B1(n1973), .Y(n2089) );
  OAI22X1 U10400 ( .A0(n199), .A1(n1974), .B0(n532), .B1(n1973), .Y(n2128) );
  OAI22X1 U10401 ( .A0(n9340), .A1(n366), .B0(n368), .B1(n2290), .Y(n2288) );
  OAI22X1 U10402 ( .A0(n9340), .A1(n186), .B0(n492), .B1(n2290), .Y(n2411) );
  NAND3X2 U10403 ( .A(N1656), .B(N1657), .C(n2132), .Y(n199) );
  MX4X1 U10404 ( .A(n9004), .B(n8994), .C(n8999), .D(n8989), .S0(n9136), .S1(
        n9137), .Y(N7386) );
  MX4X1 U10405 ( .A(n8993), .B(n8991), .C(n8992), .D(n8990), .S0(n9139), .S1(
        n9140), .Y(n8994) );
  MX4X1 U10406 ( .A(n9003), .B(n9001), .C(n9002), .D(n9000), .S0(n9139), .S1(
        n9140), .Y(n9004) );
  MX4X1 U10407 ( .A(n8988), .B(n8986), .C(n8987), .D(n8985), .S0(n9139), .S1(
        n9140), .Y(n8989) );
  CLKMX2X2 U10408 ( .A(n8530), .B(n8440), .S0(n8919), .Y(n8434) );
  CLKMX2X2 U10409 ( .A(n8550), .B(n8441), .S0(n8919), .Y(n8435) );
  NAND2X1 U10410 ( .A(avg_reg[5]), .B(n9348), .Y(n259) );
  NAND2X1 U10411 ( .A(avg_reg[6]), .B(n9348), .Y(n266) );
  NAND2X1 U10412 ( .A(avg_reg[7]), .B(n9348), .Y(n273) );
  NAND2X1 U10413 ( .A(avg_reg[9]), .B(n9348), .Y(n287) );
  MXI4X1 U10414 ( .A(n8911), .B(n8421), .C(n8743), .D(n8739), .S0(n9127), .S1(
        n8929), .Y(n8794) );
  MXI2X1 U10415 ( .A(n8740), .B(n8741), .S0(n9513), .Y(n8739) );
  CLKINVX1 U10416 ( .A(n8493), .Y(n8911) );
  MX4X1 U10417 ( .A(n8656), .B(n8650), .C(n8653), .D(n8647), .S0(n8929), .S1(
        n8926), .Y(n8659) );
  MXI2X1 U10418 ( .A(n8657), .B(n8658), .S0(n8963), .Y(n8656) );
  MX4X1 U10419 ( .A(n8669), .B(n8663), .C(n8666), .D(n8660), .S0(n8929), .S1(
        n8926), .Y(n8672) );
  MXI2X1 U10420 ( .A(n8670), .B(n8671), .S0(n8963), .Y(n8669) );
  MX4X1 U10421 ( .A(n8682), .B(n8676), .C(n8679), .D(n8673), .S0(n8929), .S1(
        n8926), .Y(n8685) );
  MXI2X1 U10422 ( .A(n8683), .B(n8684), .S0(n8963), .Y(n8682) );
  MX4X1 U10423 ( .A(n8643), .B(n8637), .C(n8640), .D(n8634), .S0(n8929), .S1(
        n8926), .Y(n8646) );
  MXI2X1 U10424 ( .A(n8644), .B(n8645), .S0(n8962), .Y(n8643) );
  MXI2X1 U10425 ( .A(n8747), .B(n8748), .S0(n9513), .Y(n8746) );
  CLKINVX1 U10426 ( .A(n8513), .Y(n8912) );
  MXI2X1 U10427 ( .A(n8754), .B(n8755), .S0(n9137), .Y(n8753) );
  CLKINVX1 U10428 ( .A(n8533), .Y(n8913) );
  CLKBUFX3 U10429 ( .A(n618), .Y(n9423) );
  OA22X1 U10430 ( .A0(n663), .A1(n230), .B0(n299), .B1(n365), .Y(n618) );
  NOR2X1 U10431 ( .A(n9780), .B(n9422), .Y(n663) );
  CLKBUFX3 U10432 ( .A(n1263), .Y(n9403) );
  OA22X1 U10433 ( .A0(n1300), .A1(n230), .B0(n299), .B1(n1024), .Y(n1263) );
  NOR2X1 U10434 ( .A(n9788), .B(n9402), .Y(n1300) );
  CLKBUFX3 U10435 ( .A(n1895), .Y(n9383) );
  OA22X1 U10436 ( .A0(n1932), .A1(n230), .B0(n299), .B1(n8187), .Y(n1895) );
  NOR2X1 U10437 ( .A(n9773), .B(n1903), .Y(n1932) );
  CLKBUFX3 U10438 ( .A(n2214), .Y(n9375) );
  OA22X1 U10439 ( .A0(n2251), .A1(n230), .B0(n299), .B1(n1974), .Y(n2214) );
  NOR2BX1 U10440 ( .AN(n9372), .B(n9374), .Y(n2251) );
  MXI4X1 U10441 ( .A(n8486), .B(n8482), .C(n8484), .D(n8480), .S0(n8927), .S1(
        n8922), .Y(n8493) );
  MXI2X1 U10442 ( .A(n8879), .B(n8487), .S0(n8963), .Y(n8486) );
  MXI3X1 U10443 ( .A(n8839), .B(n8831), .C(n8485), .S0(n8941), .S1(n8957), .Y(
        n8484) );
  MXI3X1 U10444 ( .A(n8807), .B(n8799), .C(n8481), .S0(n8941), .S1(n8957), .Y(
        n8480) );
  MXI4X1 U10445 ( .A(n8506), .B(n8502), .C(n8504), .D(n8500), .S0(n8927), .S1(
        n8922), .Y(n8513) );
  MXI2X1 U10446 ( .A(n8880), .B(n8507), .S0(n8963), .Y(n8506) );
  MXI3X1 U10447 ( .A(n8840), .B(n8832), .C(n8505), .S0(n8942), .S1(n8958), .Y(
        n8504) );
  MXI3X1 U10448 ( .A(n8808), .B(n8800), .C(n8501), .S0(n8942), .S1(n8958), .Y(
        n8500) );
  MXI4X1 U10449 ( .A(n8526), .B(n8522), .C(n8524), .D(n8520), .S0(n8927), .S1(
        n8922), .Y(n8533) );
  MXI2X1 U10450 ( .A(n8881), .B(n8527), .S0(n8963), .Y(n8526) );
  MXI3X1 U10451 ( .A(n8841), .B(n8833), .C(n8525), .S0(n8942), .S1(n8958), .Y(
        n8524) );
  MXI3X1 U10452 ( .A(n8809), .B(n8801), .C(n8521), .S0(n8942), .S1(n8958), .Y(
        n8520) );
  CLKBUFX3 U10453 ( .A(n126), .Y(n9457) );
  OA21XL U10454 ( .A0(n144), .A1(n145), .B0(n146), .Y(n126) );
  NAND4X1 U10455 ( .A(n91), .B(N1677), .C(n9744), .D(n9459), .Y(n146) );
  CLKBUFX3 U10456 ( .A(n162), .Y(n9455) );
  OA22X1 U10457 ( .A0(n159), .A1(n8263), .B0(n174), .B1(n145), .Y(n162) );
  CLKBUFX3 U10458 ( .A(n201), .Y(n9452) );
  OA22X1 U10459 ( .A0(n159), .A1(n8312), .B0(n213), .B1(n145), .Y(n201) );
  CLKBUFX3 U10460 ( .A(n214), .Y(n9451) );
  OA22X1 U10461 ( .A0(n159), .A1(n8329), .B0(n228), .B1(n145), .Y(n214) );
  CLKBUFX3 U10462 ( .A(n1580), .Y(n9393) );
  OA22X1 U10463 ( .A0(n1617), .A1(n230), .B0(n299), .B1(n1339), .Y(n1580) );
  NOR2BX1 U10464 ( .AN(n9523), .B(n9392), .Y(n1617) );
  CLKBUFX3 U10465 ( .A(n231), .Y(n9432) );
  OA22X1 U10466 ( .A0(n298), .A1(n230), .B0(n159), .B1(n299), .Y(n231) );
  NOR2X1 U10467 ( .A(n9755), .B(n9431), .Y(n298) );
  CLKBUFX3 U10468 ( .A(n175), .Y(n9454) );
  MX3XL U10469 ( .A(n8466), .B(n8905), .C(n8423), .S0(n9513), .S1(n8928), .Y(
        n8440) );
  MX3XL U10470 ( .A(n8467), .B(n8906), .C(n8424), .S0(n9137), .S1(n8928), .Y(
        n8441) );
  CLKBUFX3 U10471 ( .A(n8953), .Y(n8930) );
  CLKBUFX3 U10472 ( .A(n9509), .Y(n8953) );
  NOR2X2 U10473 ( .A(n9397), .B(n9665), .Y(n1426) );
  NOR2X2 U10474 ( .A(n9360), .B(n9665), .Y(n2420) );
  MX4X1 U10475 ( .A(n9024), .B(n9014), .C(n9019), .D(n9009), .S0(n9136), .S1(
        n9137), .Y(N7385) );
  MX4X1 U10476 ( .A(n9013), .B(n9011), .C(n9012), .D(n9010), .S0(n9139), .S1(
        n9141), .Y(n9014) );
  MX4X1 U10477 ( .A(n9023), .B(n9021), .C(n9022), .D(n9020), .S0(n9139), .S1(
        n9141), .Y(n9024) );
  MX4X1 U10478 ( .A(n9008), .B(n9006), .C(n9007), .D(n9005), .S0(n9139), .S1(
        n8431), .Y(n9009) );
  MX4X1 U10479 ( .A(n9044), .B(n9034), .C(n9039), .D(n9029), .S0(n9136), .S1(
        n9137), .Y(N7384) );
  MX4X1 U10480 ( .A(n9033), .B(n9031), .C(n9032), .D(n9030), .S0(n9138), .S1(
        n9141), .Y(n9034) );
  MX4X1 U10481 ( .A(n9043), .B(n9041), .C(n9042), .D(n9040), .S0(n9138), .S1(
        n9141), .Y(n9044) );
  MX4X1 U10482 ( .A(n9028), .B(n9026), .C(n9027), .D(n9025), .S0(n9139), .S1(
        n9141), .Y(n9029) );
  MX4X1 U10483 ( .A(n9064), .B(n9054), .C(n9059), .D(n9049), .S0(n9136), .S1(
        n9137), .Y(N7383) );
  MX4X1 U10484 ( .A(n9063), .B(n9061), .C(n9062), .D(n9060), .S0(n8928), .S1(
        n8950), .Y(n9064) );
  MX4X1 U10485 ( .A(n9053), .B(n9051), .C(n9052), .D(n9050), .S0(n8370), .S1(
        n9141), .Y(n9054) );
  MX4X1 U10486 ( .A(n9048), .B(n9046), .C(n9047), .D(n9045), .S0(n8370), .S1(
        n8940), .Y(n9049) );
  MX4X1 U10487 ( .A(n9084), .B(n9074), .C(n9079), .D(n9069), .S0(n9136), .S1(
        n9137), .Y(N7382) );
  MX4X1 U10488 ( .A(n9073), .B(n9071), .C(n9072), .D(n9070), .S0(n8370), .S1(
        n8943), .Y(n9074) );
  MX4X1 U10489 ( .A(n9083), .B(n9081), .C(n9082), .D(n9080), .S0(n8370), .S1(
        n8431), .Y(n9084) );
  MX4X1 U10490 ( .A(n9068), .B(n9066), .C(n9067), .D(n9065), .S0(n8370), .S1(
        n8431), .Y(n9069) );
  CLKMX2X2 U10491 ( .A(n8570), .B(n8446), .S0(n8919), .Y(n8442) );
  CLKMX2X2 U10492 ( .A(n8590), .B(n8447), .S0(n8919), .Y(n8443) );
  CLKMX2X2 U10493 ( .A(n8610), .B(n8448), .S0(n8919), .Y(n8444) );
  CLKMX2X2 U10494 ( .A(n8630), .B(n8449), .S0(n8919), .Y(n8445) );
  NAND2X1 U10495 ( .A(avg_reg[2]), .B(n9348), .Y(n235) );
  NAND2X1 U10496 ( .A(avg_reg[3]), .B(n9348), .Y(n245) );
  NAND2X1 U10497 ( .A(avg_reg[4]), .B(n9348), .Y(n252) );
  MX4X1 U10498 ( .A(n8695), .B(n8689), .C(n8692), .D(n8686), .S0(n8929), .S1(
        n8926), .Y(n8698) );
  MXI2X1 U10499 ( .A(n8696), .B(n8697), .S0(n8963), .Y(n8695) );
  MX4X1 U10500 ( .A(n8708), .B(n8702), .C(n8705), .D(n8699), .S0(n8929), .S1(
        n8926), .Y(n8711) );
  MXI2X1 U10501 ( .A(n8709), .B(n8710), .S0(n8962), .Y(n8708) );
  MX4X1 U10502 ( .A(n8721), .B(n8715), .C(n8718), .D(n8712), .S0(n8929), .S1(
        n8926), .Y(n8724) );
  MXI2X1 U10503 ( .A(n8722), .B(n8723), .S0(n8962), .Y(n8721) );
  MX4X1 U10504 ( .A(n8734), .B(n8728), .C(n8731), .D(n8725), .S0(n8929), .S1(
        n8926), .Y(n8737) );
  MXI2X1 U10505 ( .A(n8735), .B(n8736), .S0(n8963), .Y(n8734) );
  CLKINVX1 U10506 ( .A(n8795), .Y(N7391) );
  MXI4X1 U10507 ( .A(n8914), .B(n8424), .C(n8764), .D(n8760), .S0(n9128), .S1(
        n8929), .Y(n8795) );
  MXI2X1 U10508 ( .A(n8761), .B(n8762), .S0(n9137), .Y(n8760) );
  CLKINVX1 U10509 ( .A(n8553), .Y(n8914) );
  CLKINVX1 U10510 ( .A(n8796), .Y(N7392) );
  MXI4X1 U10511 ( .A(n8915), .B(n8426), .C(n8771), .D(n8767), .S0(n9127), .S1(
        n8929), .Y(n8796) );
  MXI2X1 U10512 ( .A(n8768), .B(n8769), .S0(n9137), .Y(n8767) );
  CLKINVX1 U10513 ( .A(n8573), .Y(n8915) );
  CLKINVX1 U10514 ( .A(n8797), .Y(N7393) );
  MXI4X1 U10515 ( .A(n8916), .B(n8425), .C(n8778), .D(n8774), .S0(n9125), .S1(
        n8929), .Y(n8797) );
  MXI2X1 U10516 ( .A(n8775), .B(n8776), .S0(n9137), .Y(n8774) );
  CLKINVX1 U10517 ( .A(n8593), .Y(n8916) );
  MXI2X1 U10518 ( .A(n8782), .B(n8783), .S0(n9137), .Y(n8781) );
  CLKINVX1 U10519 ( .A(n8613), .Y(n8917) );
  CLKINVX1 U10520 ( .A(n8798), .Y(N7395) );
  MXI4X1 U10521 ( .A(n8918), .B(n8428), .C(n8792), .D(n8788), .S0(n9127), .S1(
        n8929), .Y(n8798) );
  MXI2X1 U10522 ( .A(n8789), .B(n8790), .S0(n9137), .Y(n8788) );
  CLKINVX1 U10523 ( .A(n8633), .Y(n8918) );
  CLKBUFX3 U10524 ( .A(n1934), .Y(n9382) );
  NAND2X1 U10525 ( .A(n9459), .B(n1972), .Y(n1934) );
  OAI33X1 U10526 ( .A0(n1973), .A1(n144), .A2(n9741), .B0(n1974), .B1(n1975), 
        .B2(n982), .Y(n1972) );
  CLKBUFX3 U10527 ( .A(n943), .Y(n9413) );
  NAND2X1 U10528 ( .A(n9459), .B(n980), .Y(n943) );
  OAI31XL U10529 ( .A0(n704), .A1(n981), .A2(n982), .B0(n983), .Y(n980) );
  OAI211X1 U10530 ( .A0(n9761), .A1(n9412), .B0(n9349), .C0(n985), .Y(n983) );
  MXI4X1 U10531 ( .A(n8546), .B(n8542), .C(n8544), .D(n8540), .S0(n8927), .S1(
        n8922), .Y(n8553) );
  MXI2X1 U10532 ( .A(n8882), .B(n8547), .S0(n8963), .Y(n8546) );
  MXI3X1 U10533 ( .A(n8842), .B(n8834), .C(n8545), .S0(n8938), .S1(n8958), .Y(
        n8544) );
  MXI3X1 U10534 ( .A(n8810), .B(n8802), .C(n8541), .S0(n8945), .S1(n8958), .Y(
        n8540) );
  MXI4X1 U10535 ( .A(n8566), .B(n8562), .C(n8564), .D(n8560), .S0(n8926), .S1(
        n8923), .Y(n8573) );
  MXI2X1 U10536 ( .A(n8883), .B(n8567), .S0(n8963), .Y(n8566) );
  MXI3X1 U10537 ( .A(n8843), .B(n8835), .C(n8565), .S0(n8944), .S1(n8958), .Y(
        n8564) );
  MXI3X1 U10538 ( .A(n8811), .B(n8803), .C(n8561), .S0(n8943), .S1(n8958), .Y(
        n8560) );
  MXI4X1 U10539 ( .A(n8586), .B(n8582), .C(n8584), .D(n8580), .S0(n8927), .S1(
        n8923), .Y(n8593) );
  MXI2X1 U10540 ( .A(n8884), .B(n8587), .S0(n8963), .Y(n8586) );
  MXI3X1 U10541 ( .A(n8844), .B(n8836), .C(n8585), .S0(n8939), .S1(n8959), .Y(
        n8584) );
  MXI3X1 U10542 ( .A(n8812), .B(n8804), .C(n8581), .S0(n8940), .S1(n8958), .Y(
        n8580) );
  MXI4X1 U10543 ( .A(n8606), .B(n8602), .C(n8604), .D(n8600), .S0(n8927), .S1(
        n8922), .Y(n8613) );
  MXI2X1 U10544 ( .A(n8885), .B(n8607), .S0(n8962), .Y(n8606) );
  MXI3X1 U10545 ( .A(n8845), .B(n8837), .C(n8605), .S0(n8948), .S1(n8958), .Y(
        n8604) );
  MXI3X1 U10546 ( .A(n8813), .B(n8805), .C(n8601), .S0(n8938), .S1(n8959), .Y(
        n8600) );
  MXI4X1 U10547 ( .A(n8626), .B(n8622), .C(n8624), .D(n8620), .S0(n8926), .S1(
        n8923), .Y(n8633) );
  MXI2X1 U10548 ( .A(n8886), .B(n8627), .S0(n8963), .Y(n8626) );
  MXI3X1 U10549 ( .A(n8846), .B(n8838), .C(n8625), .S0(n8942), .S1(n8959), .Y(
        n8624) );
  MXI3X1 U10550 ( .A(n8814), .B(n8806), .C(n8621), .S0(n8946), .S1(n8959), .Y(
        n8620) );
  MX3XL U10551 ( .A(n8468), .B(n8907), .C(n8426), .S0(n8924), .S1(n8928), .Y(
        n8446) );
  MX3XL U10552 ( .A(n8469), .B(n8908), .C(n8425), .S0(n8924), .S1(n8928), .Y(
        n8447) );
  MX3XL U10553 ( .A(n8470), .B(n8909), .C(n8427), .S0(n8924), .S1(n8928), .Y(
        n8448) );
  MX3XL U10554 ( .A(n8473), .B(n8910), .C(n8428), .S0(n8925), .S1(n8928), .Y(
        n8449) );
  CLKBUFX3 U10555 ( .A(n9141), .Y(n9140) );
  CLKBUFX3 U10556 ( .A(n281), .Y(n9624) );
  CLKBUFX3 U10557 ( .A(n246), .Y(n9648) );
  CLKBUFX3 U10558 ( .A(n253), .Y(n9642) );
  CLKBUFX3 U10559 ( .A(n260), .Y(n9639) );
  MX4X1 U10560 ( .A(n9104), .B(n9094), .C(n9099), .D(n9089), .S0(n9136), .S1(
        n9137), .Y(N7381) );
  MX4X1 U10561 ( .A(n9093), .B(n9091), .C(n9092), .D(n9090), .S0(n8370), .S1(
        n8431), .Y(n9094) );
  MX4X1 U10562 ( .A(n9103), .B(n9101), .C(n9102), .D(n9100), .S0(n9511), .S1(
        n8431), .Y(n9104) );
  MX4X1 U10563 ( .A(n9088), .B(n9086), .C(n9087), .D(n9085), .S0(n8370), .S1(
        n8943), .Y(n9089) );
  MX4X1 U10564 ( .A(n9124), .B(n9114), .C(n9119), .D(n9109), .S0(n9136), .S1(
        n9137), .Y(N7380) );
  MX4X1 U10565 ( .A(n9113), .B(n9111), .C(n9112), .D(n9110), .S0(n8370), .S1(
        n8431), .Y(n9114) );
  MX4X1 U10566 ( .A(n9123), .B(n9121), .C(n9122), .D(n9120), .S0(n9511), .S1(
        n8431), .Y(n9124) );
  MX4X1 U10567 ( .A(n9108), .B(n9106), .C(n9107), .D(n9105), .S0(n9511), .S1(
        n8431), .Y(n9109) );
  NAND2X1 U10568 ( .A(IRB_RW), .B(n9339), .Y(n2565) );
  NOR2X1 U10569 ( .A(n9509), .B(n9508), .Y(n2536) );
  CLKINVX1 U10570 ( .A(n985), .Y(n9741) );
  AND2X2 U10571 ( .A(n2536), .B(n9517), .Y(n617) );
  CLKINVX1 U10572 ( .A(n9342), .Y(n9813) );
  CLKBUFX3 U10573 ( .A(n129), .Y(n9430) );
  NAND2X1 U10574 ( .A(n9341), .B(n9343), .Y(n129) );
  CLKBUFX3 U10575 ( .A(n614), .Y(n9349) );
  NAND3BX1 U10576 ( .AN(n9348), .B(n9612), .C(n9614), .Y(n614) );
  CLKBUFX3 U10577 ( .A(n292), .Y(n9613) );
  CLKBUFX3 U10578 ( .A(n94), .Y(n9660) );
  AOI221X1 U10579 ( .A0(n8370), .A1(n2546), .B0(n9510), .B1(n2541), .C0(n2538), 
        .Y(n2540) );
  AOI2BB2X1 U10580 ( .B0(n8370), .B1(n2541), .A0N(n9739), .A1N(n8370), .Y(
        n2539) );
  NAND3X2 U10581 ( .A(n8393), .B(N1661), .C(N1659), .Y(n159) );
  OAI31XL U10582 ( .A0(n9736), .A1(n2552), .A2(n9508), .B0(n9509), .Y(n2555)
         );
  CLKINVX1 U10583 ( .A(n2551), .Y(n9736) );
  OAI31XL U10584 ( .A0(n2538), .A1(n9782), .A2(n9735), .B0(n2544), .Y(n3108)
         );
  OAI31XL U10585 ( .A0(n9734), .A1(n2541), .A2(n9513), .B0(n9515), .Y(n2544)
         );
  CLKINVX1 U10586 ( .A(n2540), .Y(n9734) );
  NAND2X1 U10587 ( .A(n985), .B(n2558), .Y(n2549) );
  OAI22XL U10588 ( .A0(n2536), .A1(n9740), .B0(n9341), .B1(n9737), .Y(n2558)
         );
  NAND2X1 U10589 ( .A(n985), .B(n2547), .Y(n2538) );
  OAI22XL U10590 ( .A0(n2535), .A1(n9739), .B0(n9343), .B1(n9735), .Y(n2547)
         );
  NOR2X1 U10591 ( .A(n9515), .B(n9513), .Y(n2535) );
  NOR2X1 U10592 ( .A(n9368), .B(n9341), .Y(n144) );
  NOR2X1 U10593 ( .A(n9357), .B(n9342), .Y(n200) );
  NOR2X1 U10594 ( .A(n9362), .B(n9342), .Y(n187) );
  NAND3X1 U10595 ( .A(N1657), .B(N1658), .C(N1656), .Y(n1975) );
  BUFX4 U10596 ( .A(n676), .Y(n9410) );
  NAND2X1 U10597 ( .A(n9401), .B(n9341), .Y(n676) );
  BUFX4 U10598 ( .A(n996), .Y(n9400) );
  NAND2X1 U10599 ( .A(n9391), .B(n9341), .Y(n996) );
  BUFX4 U10600 ( .A(n1311), .Y(n9390) );
  NAND2X1 U10601 ( .A(n9344), .B(n9341), .Y(n1311) );
  BUFX4 U10602 ( .A(n1940), .Y(n9371) );
  NAND2X1 U10603 ( .A(n2211), .B(n9341), .Y(n1940) );
  BUFX4 U10604 ( .A(n2144), .Y(n9358) );
  NAND2X1 U10605 ( .A(n2211), .B(n9357), .Y(n2144) );
  BUFX4 U10606 ( .A(n384), .Y(n9419) );
  NAND2X1 U10607 ( .A(n9411), .B(n9368), .Y(n384) );
  BUFX4 U10608 ( .A(n424), .Y(n9418) );
  NAND2X1 U10609 ( .A(n9411), .B(n9365), .Y(n424) );
  BUFX4 U10610 ( .A(n464), .Y(n9417) );
  NAND2X1 U10611 ( .A(n9411), .B(n9362), .Y(n464) );
  BUFX4 U10612 ( .A(n504), .Y(n9416) );
  NAND2X1 U10613 ( .A(n9411), .B(n9342), .Y(n504) );
  BUFX4 U10614 ( .A(n544), .Y(n9415) );
  NAND2X1 U10615 ( .A(n9411), .B(n9357), .Y(n544) );
  BUFX4 U10616 ( .A(n717), .Y(n9409) );
  NAND2X1 U10617 ( .A(n9401), .B(n9368), .Y(n717) );
  BUFX4 U10618 ( .A(n756), .Y(n9408) );
  NAND2X1 U10619 ( .A(n9401), .B(n9365), .Y(n756) );
  BUFX4 U10620 ( .A(n795), .Y(n9407) );
  NAND2X1 U10621 ( .A(n9401), .B(n9362), .Y(n795) );
  BUFX4 U10622 ( .A(n834), .Y(n9406) );
  NAND2X1 U10623 ( .A(n9401), .B(n9342), .Y(n834) );
  BUFX4 U10624 ( .A(n873), .Y(n9405) );
  NAND2X1 U10625 ( .A(n9401), .B(n9357), .Y(n873) );
  BUFX4 U10626 ( .A(n1037), .Y(n9399) );
  NAND2X1 U10627 ( .A(n9391), .B(n9368), .Y(n1037) );
  BUFX4 U10628 ( .A(n1076), .Y(n9398) );
  NAND2X1 U10629 ( .A(n9391), .B(n9365), .Y(n1076) );
  BUFX4 U10630 ( .A(n1154), .Y(n9396) );
  NAND2X1 U10631 ( .A(n9391), .B(n9342), .Y(n1154) );
  BUFX4 U10632 ( .A(n1193), .Y(n9395) );
  NAND2X1 U10633 ( .A(n9391), .B(n9357), .Y(n1193) );
  BUFX4 U10634 ( .A(n1352), .Y(n9389) );
  NAND2X1 U10635 ( .A(n9344), .B(n9368), .Y(n1352) );
  BUFX4 U10636 ( .A(n1427), .Y(n9387) );
  NAND2X1 U10637 ( .A(n9344), .B(n9362), .Y(n1427) );
  BUFX4 U10638 ( .A(n1510), .Y(n9385) );
  NAND2X1 U10639 ( .A(n9344), .B(n9357), .Y(n1510) );
  BUFX4 U10640 ( .A(n1667), .Y(n9381) );
  NAND2X1 U10641 ( .A(n9373), .B(n9368), .Y(n1667) );
  BUFX4 U10642 ( .A(n1706), .Y(n9380) );
  NAND2X1 U10643 ( .A(n9373), .B(n9365), .Y(n1706) );
  BUFX4 U10644 ( .A(n1745), .Y(n9379) );
  NAND2X1 U10645 ( .A(n9373), .B(n9362), .Y(n1745) );
  BUFX4 U10646 ( .A(n1784), .Y(n9378) );
  NAND2X1 U10647 ( .A(n9373), .B(n9342), .Y(n1784) );
  BUFX4 U10648 ( .A(n1825), .Y(n9377) );
  NAND2X1 U10649 ( .A(n9373), .B(n9357), .Y(n1825) );
  NAND2X1 U10650 ( .A(n9411), .B(n9341), .Y(n312) );
  BUFX4 U10651 ( .A(n1391), .Y(n9388) );
  NAND2X1 U10652 ( .A(n9344), .B(n9365), .Y(n1391) );
  NOR3X1 U10653 ( .A(n9510), .B(n9512), .C(n9515), .Y(n1577) );
  BUFX4 U10654 ( .A(n1984), .Y(n9369) );
  NAND2X1 U10655 ( .A(n2211), .B(n9368), .Y(n1984) );
  BUFX4 U10656 ( .A(n2023), .Y(n9366) );
  NAND2X1 U10657 ( .A(n2211), .B(n9365), .Y(n2023) );
  BUFX4 U10658 ( .A(n2062), .Y(n9363) );
  NAND2X1 U10659 ( .A(n2211), .B(n9362), .Y(n2062) );
  NAND2X1 U10660 ( .A(n9368), .B(n9343), .Y(n151) );
  NAND2X1 U10661 ( .A(n9365), .B(n9343), .Y(n165) );
  NAND2X1 U10662 ( .A(n9362), .B(n9343), .Y(n178) );
  NAND2X1 U10663 ( .A(n9342), .B(n9343), .Y(n191) );
  NAND2X1 U10664 ( .A(n9357), .B(n9343), .Y(n204) );
  INVX3 U10665 ( .A(n9339), .Y(n9744) );
  CLKINVX1 U10666 ( .A(n2552), .Y(n9737) );
  CLKINVX1 U10667 ( .A(n2541), .Y(n9735) );
  NOR2X1 U10668 ( .A(n9357), .B(n617), .Y(n213) );
  NOR2X1 U10669 ( .A(n9368), .B(n9365), .Y(n161) );
  NOR2X1 U10670 ( .A(n9365), .B(n9362), .Y(n174) );
  CLKINVX1 U10671 ( .A(n91), .Y(n9746) );
  NOR3X1 U10672 ( .A(n9510), .B(n9514), .C(n9513), .Y(n940) );
  CLKBUFX3 U10673 ( .A(n1260), .Y(n9391) );
  CLKBUFX3 U10674 ( .A(n1892), .Y(n9373) );
  CLKINVX1 U10675 ( .A(n2546), .Y(n9739) );
  CLKINVX1 U10676 ( .A(n2557), .Y(n9740) );
  CLKBUFX3 U10677 ( .A(n2252), .Y(n9372) );
  NAND2X1 U10678 ( .A(n2294), .B(n9341), .Y(n2252) );
  CLKBUFX3 U10679 ( .A(n2421), .Y(n9361) );
  NAND2X1 U10680 ( .A(n2294), .B(n9342), .Y(n2421) );
  CLKBUFX3 U10681 ( .A(n2303), .Y(n9370) );
  NAND2X1 U10682 ( .A(n2294), .B(n9368), .Y(n2303) );
  CLKBUFX3 U10683 ( .A(n2343), .Y(n9367) );
  NAND2X1 U10684 ( .A(n2294), .B(n9365), .Y(n2343) );
  CLKBUFX3 U10685 ( .A(n2383), .Y(n9364) );
  NAND2X1 U10686 ( .A(n2294), .B(n9362), .Y(n2383) );
  CLKBUFX3 U10687 ( .A(n2462), .Y(n9359) );
  NAND2X1 U10688 ( .A(n2294), .B(n9357), .Y(n2462) );
  AND2X2 U10689 ( .A(n2535), .B(n9511), .Y(n2211) );
  CLKINVX1 U10690 ( .A(n9606), .Y(n9612) );
  NOR3X1 U10691 ( .A(n9748), .B(n9738), .C(n9747), .Y(n92) );
  CLKINVX1 U10692 ( .A(n96), .Y(n9745) );
  MX4X1 U10693 ( .A(n9157), .B(n9155), .C(n9156), .D(n9154), .S0(n9337), .S1(
        n9333), .Y(n9158) );
  MX4X1 U10694 ( .A(n9162), .B(n9160), .C(n9161), .D(n9159), .S0(n9337), .S1(
        n9334), .Y(n9163) );
  MX4X1 U10695 ( .A(n9177), .B(n9175), .C(n9176), .D(n9174), .S0(n9337), .S1(
        n9334), .Y(n9178) );
  MX4X1 U10696 ( .A(n9187), .B(n9185), .C(n9186), .D(n9184), .S0(n9335), .S1(
        n9333), .Y(n9188) );
  MX4X1 U10697 ( .A(n9197), .B(n9195), .C(n9196), .D(n9194), .S0(n9335), .S1(
        n9333), .Y(n9198) );
  MX4X1 U10698 ( .A(n9207), .B(n9205), .C(n9206), .D(n9204), .S0(n9335), .S1(
        n9333), .Y(n9208) );
  MX4X1 U10699 ( .A(n9217), .B(n9215), .C(n9216), .D(n9214), .S0(n9335), .S1(
        n9333), .Y(n9218) );
  MX4X1 U10700 ( .A(n9227), .B(n9225), .C(n9226), .D(n9224), .S0(n9335), .S1(
        n9333), .Y(n9228) );
  MX4X1 U10701 ( .A(n9252), .B(n9250), .C(n9251), .D(n9249), .S0(n9336), .S1(
        n9334), .Y(n9253) );
  MX4X1 U10702 ( .A(n9237), .B(n9235), .C(n9236), .D(n9234), .S0(n9335), .S1(
        n9333), .Y(n9238) );
  MX4X1 U10703 ( .A(n9257), .B(n9255), .C(n9256), .D(n9254), .S0(n9336), .S1(
        n9333), .Y(n9258) );
  MX4X1 U10704 ( .A(n9267), .B(n9265), .C(n9266), .D(n9264), .S0(n9336), .S1(
        n9334), .Y(n9268) );
  MX4X1 U10705 ( .A(n9293), .B(n9283), .C(n9288), .D(n9278), .S0(N1661), .S1(
        n8393), .Y(N7372) );
  MX4X1 U10706 ( .A(n9277), .B(n9275), .C(n9276), .D(n9274), .S0(n9336), .S1(
        n9334), .Y(n9278) );
  MX4X1 U10707 ( .A(n9287), .B(n9285), .C(n9286), .D(n9284), .S0(n9336), .S1(
        n9334), .Y(n9288) );
  MX4X1 U10708 ( .A(n9313), .B(n9303), .C(n9308), .D(n9298), .S0(N1661), .S1(
        n8393), .Y(N7371) );
  MX4X1 U10709 ( .A(n9297), .B(n9295), .C(n9296), .D(n9294), .S0(n9336), .S1(
        n9334), .Y(n9298) );
  MX4X1 U10710 ( .A(n9307), .B(n9305), .C(n9306), .D(n9304), .S0(n9336), .S1(
        n9334), .Y(n9308) );
  MX4X1 U10711 ( .A(\buff[36][0] ), .B(\buff[37][0] ), .C(\buff[38][0] ), .D(
        \buff[39][0] ), .S0(n9317), .S1(n9328), .Y(n9161) );
  MX4X1 U10712 ( .A(\buff[4][4] ), .B(\buff[5][4] ), .C(\buff[6][4] ), .D(
        \buff[7][4] ), .S0(n9323), .S1(n9328), .Y(n9251) );
  MX4X1 U10713 ( .A(n9167), .B(n9165), .C(n9166), .D(n9164), .S0(n9337), .S1(
        n9334), .Y(n9168) );
  MX4X1 U10714 ( .A(\buff[28][0] ), .B(\buff[29][0] ), .C(\buff[30][0] ), .D(
        \buff[31][0] ), .S0(n9317), .S1(n9328), .Y(n9164) );
  MX4X1 U10715 ( .A(\buff[20][0] ), .B(\buff[21][0] ), .C(\buff[22][0] ), .D(
        \buff[23][0] ), .S0(n9317), .S1(n9330), .Y(n9166) );
  MX4X1 U10716 ( .A(\buff[24][0] ), .B(\buff[25][0] ), .C(\buff[26][0] ), .D(
        \buff[27][0] ), .S0(n9317), .S1(n9331), .Y(n9165) );
  MX4X1 U10717 ( .A(\buff[20][1] ), .B(\buff[21][1] ), .C(\buff[22][1] ), .D(
        \buff[23][1] ), .S0(n9319), .S1(n9325), .Y(n9186) );
  MX4X1 U10718 ( .A(\buff[52][1] ), .B(\buff[53][1] ), .C(\buff[54][1] ), .D(
        \buff[55][1] ), .S0(n9318), .S1(n9331), .Y(n9176) );
  MX4X1 U10719 ( .A(\buff[20][2] ), .B(\buff[21][2] ), .C(\buff[22][2] ), .D(
        \buff[23][2] ), .S0(n9320), .S1(n9326), .Y(n9206) );
  MX4X1 U10720 ( .A(\buff[52][2] ), .B(\buff[53][2] ), .C(\buff[54][2] ), .D(
        \buff[55][2] ), .S0(n9319), .S1(n9325), .Y(n9196) );
  MX4X1 U10721 ( .A(\buff[20][3] ), .B(\buff[21][3] ), .C(\buff[22][3] ), .D(
        \buff[23][3] ), .S0(n9321), .S1(n9327), .Y(n9226) );
  MX4X1 U10722 ( .A(\buff[52][3] ), .B(\buff[53][3] ), .C(\buff[54][3] ), .D(
        \buff[55][3] ), .S0(n9321), .S1(n9327), .Y(n9216) );
  MX4X1 U10723 ( .A(\buff[52][4] ), .B(\buff[53][4] ), .C(\buff[54][4] ), .D(
        \buff[55][4] ), .S0(n9322), .S1(n9327), .Y(n9236) );
  MX4X1 U10724 ( .A(\buff[20][5] ), .B(\buff[21][5] ), .C(\buff[22][5] ), .D(
        \buff[23][5] ), .S0(n9324), .S1(n9329), .Y(n9266) );
  MX4X1 U10725 ( .A(\buff[52][5] ), .B(\buff[53][5] ), .C(\buff[54][5] ), .D(
        \buff[55][5] ), .S0(n9323), .S1(n9328), .Y(n9256) );
  MX4X1 U10726 ( .A(\buff[20][6] ), .B(\buff[21][6] ), .C(\buff[22][6] ), .D(
        \buff[23][6] ), .S0(n9314), .S1(n9330), .Y(n9286) );
  MX4X1 U10727 ( .A(\buff[52][6] ), .B(\buff[53][6] ), .C(\buff[54][6] ), .D(
        \buff[55][6] ), .S0(n9324), .S1(n9329), .Y(n9276) );
  MX4X1 U10728 ( .A(\buff[20][7] ), .B(\buff[21][7] ), .C(\buff[22][7] ), .D(
        \buff[23][7] ), .S0(n9314), .S1(n9331), .Y(n9306) );
  MX4X1 U10729 ( .A(\buff[52][7] ), .B(\buff[53][7] ), .C(\buff[54][7] ), .D(
        \buff[55][7] ), .S0(n9315), .S1(n9330), .Y(n9296) );
  MX4X1 U10730 ( .A(n9247), .B(n9245), .C(n9246), .D(n9244), .S0(n9335), .S1(
        n9333), .Y(n9248) );
  MX4X1 U10731 ( .A(\buff[28][4] ), .B(\buff[29][4] ), .C(\buff[30][4] ), .D(
        \buff[31][4] ), .S0(n9322), .S1(n9326), .Y(n9244) );
  MX4X1 U10732 ( .A(\buff[20][4] ), .B(\buff[21][4] ), .C(\buff[22][4] ), .D(
        \buff[23][4] ), .S0(n9322), .S1(n9326), .Y(n9246) );
  MX4X1 U10733 ( .A(\buff[24][4] ), .B(\buff[25][4] ), .C(\buff[26][4] ), .D(
        \buff[27][4] ), .S0(n9322), .S1(n9327), .Y(n9245) );
  MX4X1 U10734 ( .A(\buff[52][0] ), .B(\buff[53][0] ), .C(\buff[54][0] ), .D(
        \buff[55][0] ), .S0(n9317), .S1(n9330), .Y(n9156) );
  MX4X1 U10735 ( .A(\buff[0][0] ), .B(\buff[1][0] ), .C(\buff[2][0] ), .D(
        \buff[3][0] ), .S0(n9318), .S1(n9332), .Y(n9172) );
  MX4X1 U10736 ( .A(\buff[16][0] ), .B(\buff[17][0] ), .C(\buff[18][0] ), .D(
        \buff[19][0] ), .S0(n9318), .S1(n9331), .Y(n9167) );
  MX4X1 U10737 ( .A(\buff[32][0] ), .B(\buff[33][0] ), .C(\buff[34][0] ), .D(
        \buff[35][0] ), .S0(n9317), .S1(N1657), .Y(n9162) );
  MX4X1 U10738 ( .A(\buff[48][0] ), .B(\buff[49][0] ), .C(\buff[50][0] ), .D(
        \buff[51][0] ), .S0(n9317), .S1(n9330), .Y(n9157) );
  MX4X1 U10739 ( .A(\buff[0][1] ), .B(\buff[1][1] ), .C(\buff[2][1] ), .D(
        \buff[3][1] ), .S0(n9319), .S1(n9325), .Y(n9192) );
  MX4X1 U10740 ( .A(\buff[32][1] ), .B(\buff[33][1] ), .C(\buff[34][1] ), .D(
        \buff[35][1] ), .S0(n9318), .S1(n9332), .Y(n9182) );
  MX4X1 U10741 ( .A(\buff[16][1] ), .B(\buff[17][1] ), .C(\buff[18][1] ), .D(
        \buff[19][1] ), .S0(n9319), .S1(n9325), .Y(n9187) );
  MX4X1 U10742 ( .A(\buff[48][1] ), .B(\buff[49][1] ), .C(\buff[50][1] ), .D(
        \buff[51][1] ), .S0(n9318), .S1(n9331), .Y(n9177) );
  MX4X1 U10743 ( .A(\buff[0][2] ), .B(\buff[1][2] ), .C(\buff[2][2] ), .D(
        \buff[3][2] ), .S0(n9320), .S1(n9326), .Y(n9212) );
  MX4X1 U10744 ( .A(\buff[32][2] ), .B(\buff[33][2] ), .C(\buff[34][2] ), .D(
        \buff[35][2] ), .S0(n9320), .S1(n9326), .Y(n9202) );
  MX4X1 U10745 ( .A(\buff[16][2] ), .B(\buff[17][2] ), .C(\buff[18][2] ), .D(
        \buff[19][2] ), .S0(n9320), .S1(n9326), .Y(n9207) );
  MX4X1 U10746 ( .A(\buff[48][2] ), .B(\buff[49][2] ), .C(\buff[50][2] ), .D(
        \buff[51][2] ), .S0(n9319), .S1(n9325), .Y(n9197) );
  MX4X1 U10747 ( .A(\buff[0][3] ), .B(\buff[1][3] ), .C(\buff[2][3] ), .D(
        \buff[3][3] ), .S0(n9322), .S1(n9326), .Y(n9232) );
  MX4X1 U10748 ( .A(\buff[32][3] ), .B(\buff[33][3] ), .C(\buff[34][3] ), .D(
        \buff[35][3] ), .S0(n9321), .S1(n9327), .Y(n9222) );
  MX4X1 U10749 ( .A(\buff[16][3] ), .B(\buff[17][3] ), .C(\buff[18][3] ), .D(
        \buff[19][3] ), .S0(n9321), .S1(n9327), .Y(n9227) );
  MX4X1 U10750 ( .A(\buff[48][3] ), .B(\buff[49][3] ), .C(\buff[50][3] ), .D(
        \buff[51][3] ), .S0(n9321), .S1(n9327), .Y(n9217) );
  MX4X1 U10751 ( .A(\buff[32][4] ), .B(\buff[33][4] ), .C(\buff[34][4] ), .D(
        \buff[35][4] ), .S0(n9322), .S1(n9327), .Y(n9242) );
  MX4X1 U10752 ( .A(\buff[16][4] ), .B(\buff[17][4] ), .C(\buff[18][4] ), .D(
        \buff[19][4] ), .S0(n9322), .S1(n9327), .Y(n9247) );
  MX4X1 U10753 ( .A(\buff[48][4] ), .B(\buff[49][4] ), .C(\buff[50][4] ), .D(
        \buff[51][4] ), .S0(n9322), .S1(n9326), .Y(n9237) );
  MX4X1 U10754 ( .A(\buff[0][4] ), .B(\buff[1][4] ), .C(\buff[2][4] ), .D(
        \buff[3][4] ), .S0(n9323), .S1(n9328), .Y(n9252) );
  MX4X1 U10755 ( .A(\buff[0][5] ), .B(\buff[1][5] ), .C(\buff[2][5] ), .D(
        \buff[3][5] ), .S0(n9324), .S1(n9329), .Y(n9272) );
  MX4X1 U10756 ( .A(\buff[32][5] ), .B(\buff[33][5] ), .C(\buff[34][5] ), .D(
        \buff[35][5] ), .S0(n9323), .S1(n9328), .Y(n9262) );
  MX4X1 U10757 ( .A(\buff[16][5] ), .B(\buff[17][5] ), .C(\buff[18][5] ), .D(
        \buff[19][5] ), .S0(n9324), .S1(n9329), .Y(n9267) );
  MX4X1 U10758 ( .A(\buff[48][5] ), .B(\buff[49][5] ), .C(\buff[50][5] ), .D(
        \buff[51][5] ), .S0(n9323), .S1(n9328), .Y(n9257) );
  MX4X1 U10759 ( .A(\buff[0][6] ), .B(\buff[1][6] ), .C(\buff[2][6] ), .D(
        \buff[3][6] ), .S0(n9316), .S1(n9330), .Y(n9292) );
  MX4X1 U10760 ( .A(\buff[32][6] ), .B(\buff[33][6] ), .C(\buff[34][6] ), .D(
        \buff[35][6] ), .S0(n9314), .S1(n9330), .Y(n9282) );
  MX4X1 U10761 ( .A(\buff[16][6] ), .B(\buff[17][6] ), .C(\buff[18][6] ), .D(
        \buff[19][6] ), .S0(n9316), .S1(n9330), .Y(n9287) );
  MX4X1 U10762 ( .A(\buff[48][6] ), .B(\buff[49][6] ), .C(\buff[50][6] ), .D(
        \buff[51][6] ), .S0(n9324), .S1(n9329), .Y(n9277) );
  MX4X1 U10763 ( .A(\buff[0][7] ), .B(\buff[1][7] ), .C(\buff[2][7] ), .D(
        \buff[3][7] ), .S0(n9314), .S1(n9331), .Y(n9312) );
  MX4X1 U10764 ( .A(\buff[32][7] ), .B(\buff[33][7] ), .C(\buff[34][7] ), .D(
        \buff[35][7] ), .S0(n9315), .S1(n9331), .Y(n9302) );
  MX4X1 U10765 ( .A(\buff[16][7] ), .B(\buff[17][7] ), .C(\buff[18][7] ), .D(
        \buff[19][7] ), .S0(n9316), .S1(n9331), .Y(n9307) );
  MX4X1 U10766 ( .A(\buff[48][7] ), .B(\buff[49][7] ), .C(\buff[50][7] ), .D(
        \buff[51][7] ), .S0(n9315), .S1(n9331), .Y(n9297) );
  MX4X1 U10767 ( .A(n9172), .B(n9170), .C(n9171), .D(n9169), .S0(n9337), .S1(
        n9334), .Y(n9173) );
  MX4X1 U10768 ( .A(\buff[12][0] ), .B(\buff[13][0] ), .C(\buff[14][0] ), .D(
        \buff[15][0] ), .S0(n9318), .S1(n9332), .Y(n9169) );
  MX4X1 U10769 ( .A(\buff[4][0] ), .B(\buff[5][0] ), .C(\buff[6][0] ), .D(
        \buff[7][0] ), .S0(n9318), .S1(N1657), .Y(n9171) );
  MX4X1 U10770 ( .A(\buff[8][0] ), .B(\buff[9][0] ), .C(\buff[10][0] ), .D(
        \buff[11][0] ), .S0(n9318), .S1(n9332), .Y(n9170) );
  MX4X1 U10771 ( .A(n9192), .B(n9190), .C(n9191), .D(n9189), .S0(n9335), .S1(
        n9333), .Y(n9193) );
  MX4X1 U10772 ( .A(\buff[12][1] ), .B(\buff[13][1] ), .C(\buff[14][1] ), .D(
        \buff[15][1] ), .S0(n9319), .S1(n9325), .Y(n9189) );
  MX4X1 U10773 ( .A(\buff[4][1] ), .B(\buff[5][1] ), .C(\buff[6][1] ), .D(
        \buff[7][1] ), .S0(n9319), .S1(n9325), .Y(n9191) );
  MX4X1 U10774 ( .A(\buff[8][1] ), .B(\buff[9][1] ), .C(\buff[10][1] ), .D(
        \buff[11][1] ), .S0(n9319), .S1(n9325), .Y(n9190) );
  MX4X1 U10775 ( .A(n9212), .B(n9210), .C(n9211), .D(n9209), .S0(n9335), .S1(
        n9333), .Y(n9213) );
  MX4X1 U10776 ( .A(\buff[12][2] ), .B(\buff[13][2] ), .C(\buff[14][2] ), .D(
        \buff[15][2] ), .S0(n9320), .S1(n9326), .Y(n9209) );
  MX4X1 U10777 ( .A(\buff[4][2] ), .B(\buff[5][2] ), .C(\buff[6][2] ), .D(
        \buff[7][2] ), .S0(n9320), .S1(n9326), .Y(n9211) );
  MX4X1 U10778 ( .A(\buff[8][2] ), .B(\buff[9][2] ), .C(\buff[10][2] ), .D(
        \buff[11][2] ), .S0(n9320), .S1(n9326), .Y(n9210) );
  MX4X1 U10779 ( .A(n9232), .B(n9230), .C(n9231), .D(n9229), .S0(n9335), .S1(
        n9333), .Y(n9233) );
  MX4X1 U10780 ( .A(\buff[12][3] ), .B(\buff[13][3] ), .C(\buff[14][3] ), .D(
        \buff[15][3] ), .S0(n9321), .S1(n9327), .Y(n9229) );
  MX4X1 U10781 ( .A(\buff[4][3] ), .B(\buff[5][3] ), .C(\buff[6][3] ), .D(
        \buff[7][3] ), .S0(n9321), .S1(n9327), .Y(n9231) );
  MX4X1 U10782 ( .A(\buff[8][3] ), .B(\buff[9][3] ), .C(\buff[10][3] ), .D(
        \buff[11][3] ), .S0(n9321), .S1(n9327), .Y(n9230) );
  MX4X1 U10783 ( .A(n9272), .B(n9270), .C(n9271), .D(n9269), .S0(n9336), .S1(
        n9334), .Y(n9273) );
  MX4X1 U10784 ( .A(\buff[12][5] ), .B(\buff[13][5] ), .C(\buff[14][5] ), .D(
        \buff[15][5] ), .S0(n9324), .S1(n9329), .Y(n9269) );
  MX4X1 U10785 ( .A(\buff[4][5] ), .B(\buff[5][5] ), .C(\buff[6][5] ), .D(
        \buff[7][5] ), .S0(n9324), .S1(n9329), .Y(n9271) );
  MX4X1 U10786 ( .A(\buff[8][5] ), .B(\buff[9][5] ), .C(\buff[10][5] ), .D(
        \buff[11][5] ), .S0(n9324), .S1(n9329), .Y(n9270) );
  MX4X1 U10787 ( .A(n9292), .B(n9290), .C(n9291), .D(n9289), .S0(n9336), .S1(
        n9334), .Y(n9293) );
  MX4X1 U10788 ( .A(\buff[12][6] ), .B(\buff[13][6] ), .C(\buff[14][6] ), .D(
        \buff[15][6] ), .S0(n9315), .S1(n9330), .Y(n9289) );
  MX4X1 U10789 ( .A(\buff[4][6] ), .B(\buff[5][6] ), .C(\buff[6][6] ), .D(
        \buff[7][6] ), .S0(N1656), .S1(n9330), .Y(n9291) );
  MX4X1 U10790 ( .A(\buff[8][6] ), .B(\buff[9][6] ), .C(\buff[10][6] ), .D(
        \buff[11][6] ), .S0(n9316), .S1(n9330), .Y(n9290) );
  MX4X1 U10791 ( .A(n9312), .B(n9310), .C(n9311), .D(n9309), .S0(n9336), .S1(
        n9334), .Y(n9313) );
  MX4X1 U10792 ( .A(\buff[12][7] ), .B(\buff[13][7] ), .C(\buff[14][7] ), .D(
        \buff[15][7] ), .S0(n9316), .S1(n9331), .Y(n9309) );
  MX4X1 U10793 ( .A(\buff[4][7] ), .B(\buff[5][7] ), .C(\buff[6][7] ), .D(
        \buff[7][7] ), .S0(N1656), .S1(n9331), .Y(n9311) );
  MX4X1 U10794 ( .A(\buff[8][7] ), .B(\buff[9][7] ), .C(\buff[10][7] ), .D(
        \buff[11][7] ), .S0(n9314), .S1(n9331), .Y(n9310) );
  MX4X1 U10795 ( .A(\buff[44][0] ), .B(\buff[45][0] ), .C(\buff[46][0] ), .D(
        \buff[47][0] ), .S0(n9317), .S1(N1657), .Y(n9159) );
  MX4X1 U10796 ( .A(\buff[28][1] ), .B(\buff[29][1] ), .C(\buff[30][1] ), .D(
        \buff[31][1] ), .S0(n9319), .S1(n9325), .Y(n9184) );
  MX4X1 U10797 ( .A(\buff[28][2] ), .B(\buff[29][2] ), .C(\buff[30][2] ), .D(
        \buff[31][2] ), .S0(n9320), .S1(n9326), .Y(n9204) );
  MX4X1 U10798 ( .A(\buff[28][3] ), .B(\buff[29][3] ), .C(\buff[30][3] ), .D(
        \buff[31][3] ), .S0(n9321), .S1(n9327), .Y(n9224) );
  MX4X1 U10799 ( .A(\buff[12][4] ), .B(\buff[13][4] ), .C(\buff[14][4] ), .D(
        \buff[15][4] ), .S0(n9323), .S1(n9328), .Y(n9249) );
  MX4X1 U10800 ( .A(\buff[28][5] ), .B(\buff[29][5] ), .C(\buff[30][5] ), .D(
        \buff[31][5] ), .S0(n9323), .S1(n9328), .Y(n9264) );
  MX4X1 U10801 ( .A(\buff[28][6] ), .B(\buff[29][6] ), .C(\buff[30][6] ), .D(
        \buff[31][6] ), .S0(n9314), .S1(n9330), .Y(n9284) );
  MX4X1 U10802 ( .A(\buff[28][7] ), .B(\buff[29][7] ), .C(\buff[30][7] ), .D(
        \buff[31][7] ), .S0(n9315), .S1(n9331), .Y(n9304) );
  MX4X1 U10803 ( .A(\buff[60][1] ), .B(\buff[61][1] ), .C(\buff[62][1] ), .D(
        \buff[63][1] ), .S0(n9318), .S1(n9329), .Y(n9174) );
  MX4X1 U10804 ( .A(\buff[60][2] ), .B(\buff[61][2] ), .C(\buff[62][2] ), .D(
        \buff[63][2] ), .S0(n9319), .S1(n9325), .Y(n9194) );
  MX4X1 U10805 ( .A(\buff[60][3] ), .B(\buff[61][3] ), .C(\buff[62][3] ), .D(
        \buff[63][3] ), .S0(n9320), .S1(n9326), .Y(n9214) );
  MX4X1 U10806 ( .A(\buff[60][4] ), .B(\buff[61][4] ), .C(\buff[62][4] ), .D(
        \buff[63][4] ), .S0(n9322), .S1(n9325), .Y(n9234) );
  MX4X1 U10807 ( .A(\buff[60][5] ), .B(\buff[61][5] ), .C(\buff[62][5] ), .D(
        \buff[63][5] ), .S0(n9323), .S1(n9328), .Y(n9254) );
  MX4X1 U10808 ( .A(\buff[60][6] ), .B(\buff[61][6] ), .C(\buff[62][6] ), .D(
        \buff[63][6] ), .S0(n9324), .S1(n9329), .Y(n9274) );
  MX4X1 U10809 ( .A(\buff[60][7] ), .B(\buff[61][7] ), .C(\buff[62][7] ), .D(
        \buff[63][7] ), .S0(n9316), .S1(n9330), .Y(n9294) );
  MX4X1 U10810 ( .A(\buff[60][0] ), .B(\buff[61][0] ), .C(\buff[62][0] ), .D(
        \buff[63][0] ), .S0(n9317), .S1(n9330), .Y(n9154) );
  MX4X1 U10811 ( .A(\buff[40][0] ), .B(\buff[41][0] ), .C(\buff[42][0] ), .D(
        \buff[43][0] ), .S0(n9317), .S1(n9329), .Y(n9160) );
  MX4X1 U10812 ( .A(\buff[8][4] ), .B(\buff[9][4] ), .C(\buff[10][4] ), .D(
        \buff[11][4] ), .S0(n9323), .S1(n9328), .Y(n9250) );
  MX4X1 U10813 ( .A(n9182), .B(n9180), .C(n9181), .D(n9179), .S0(n9337), .S1(
        n9334), .Y(n9183) );
  MX4X1 U10814 ( .A(\buff[44][1] ), .B(\buff[45][1] ), .C(\buff[46][1] ), .D(
        \buff[47][1] ), .S0(n9318), .S1(n9332), .Y(n9179) );
  MX4X1 U10815 ( .A(\buff[36][1] ), .B(\buff[37][1] ), .C(\buff[38][1] ), .D(
        \buff[39][1] ), .S0(n9318), .S1(n9328), .Y(n9181) );
  MX4X1 U10816 ( .A(\buff[40][1] ), .B(\buff[41][1] ), .C(\buff[42][1] ), .D(
        \buff[43][1] ), .S0(n9318), .S1(n9332), .Y(n9180) );
  MX4X1 U10817 ( .A(\buff[24][1] ), .B(\buff[25][1] ), .C(\buff[26][1] ), .D(
        \buff[27][1] ), .S0(n9319), .S1(n9325), .Y(n9185) );
  MX4X1 U10818 ( .A(\buff[56][1] ), .B(\buff[57][1] ), .C(\buff[58][1] ), .D(
        \buff[59][1] ), .S0(n9318), .S1(n9329), .Y(n9175) );
  MX4X1 U10819 ( .A(\buff[24][2] ), .B(\buff[25][2] ), .C(\buff[26][2] ), .D(
        \buff[27][2] ), .S0(n9320), .S1(n9326), .Y(n9205) );
  MX4X1 U10820 ( .A(\buff[56][2] ), .B(\buff[57][2] ), .C(\buff[58][2] ), .D(
        \buff[59][2] ), .S0(n9319), .S1(n9325), .Y(n9195) );
  MX4X1 U10821 ( .A(\buff[24][3] ), .B(\buff[25][3] ), .C(\buff[26][3] ), .D(
        \buff[27][3] ), .S0(n9321), .S1(n9327), .Y(n9225) );
  MX4X1 U10822 ( .A(\buff[56][3] ), .B(\buff[57][3] ), .C(\buff[58][3] ), .D(
        \buff[59][3] ), .S0(n9320), .S1(n9326), .Y(n9215) );
  MX4X1 U10823 ( .A(\buff[56][4] ), .B(\buff[57][4] ), .C(\buff[58][4] ), .D(
        \buff[59][4] ), .S0(n9322), .S1(n9325), .Y(n9235) );
  MX4X1 U10824 ( .A(\buff[24][5] ), .B(\buff[25][5] ), .C(\buff[26][5] ), .D(
        \buff[27][5] ), .S0(n9324), .S1(n9329), .Y(n9265) );
  MX4X1 U10825 ( .A(\buff[56][5] ), .B(\buff[57][5] ), .C(\buff[58][5] ), .D(
        \buff[59][5] ), .S0(n9323), .S1(n9328), .Y(n9255) );
  MX4X1 U10826 ( .A(\buff[24][6] ), .B(\buff[25][6] ), .C(\buff[26][6] ), .D(
        \buff[27][6] ), .S0(n9315), .S1(n9330), .Y(n9285) );
  MX4X1 U10827 ( .A(\buff[56][6] ), .B(\buff[57][6] ), .C(\buff[58][6] ), .D(
        \buff[59][6] ), .S0(n9324), .S1(n9329), .Y(n9275) );
  MX4X1 U10828 ( .A(\buff[24][7] ), .B(\buff[25][7] ), .C(\buff[26][7] ), .D(
        \buff[27][7] ), .S0(n9316), .S1(n9331), .Y(n9305) );
  MX4X1 U10829 ( .A(\buff[56][7] ), .B(\buff[57][7] ), .C(\buff[58][7] ), .D(
        \buff[59][7] ), .S0(n9315), .S1(n9330), .Y(n9295) );
  MX4X1 U10830 ( .A(n9202), .B(n9200), .C(n9201), .D(n9199), .S0(n9335), .S1(
        n9333), .Y(n9203) );
  MX4X1 U10831 ( .A(\buff[44][2] ), .B(\buff[45][2] ), .C(\buff[46][2] ), .D(
        \buff[47][2] ), .S0(n9319), .S1(n9325), .Y(n9199) );
  MX4X1 U10832 ( .A(\buff[36][2] ), .B(\buff[37][2] ), .C(\buff[38][2] ), .D(
        \buff[39][2] ), .S0(n9320), .S1(n9326), .Y(n9201) );
  MX4X1 U10833 ( .A(\buff[40][2] ), .B(\buff[41][2] ), .C(\buff[42][2] ), .D(
        \buff[43][2] ), .S0(n9320), .S1(n9326), .Y(n9200) );
  MX4X1 U10834 ( .A(n9222), .B(n9220), .C(n9221), .D(n9219), .S0(n9335), .S1(
        n9333), .Y(n9223) );
  MX4X1 U10835 ( .A(\buff[44][3] ), .B(\buff[45][3] ), .C(\buff[46][3] ), .D(
        \buff[47][3] ), .S0(n9321), .S1(n9327), .Y(n9219) );
  MX4X1 U10836 ( .A(\buff[36][3] ), .B(\buff[37][3] ), .C(\buff[38][3] ), .D(
        \buff[39][3] ), .S0(n9321), .S1(n9327), .Y(n9221) );
  MX4X1 U10837 ( .A(\buff[40][3] ), .B(\buff[41][3] ), .C(\buff[42][3] ), .D(
        \buff[43][3] ), .S0(n9321), .S1(n9327), .Y(n9220) );
  MX4X1 U10838 ( .A(n9242), .B(n9240), .C(n9241), .D(n9239), .S0(n9335), .S1(
        n9333), .Y(n9243) );
  MX4X1 U10839 ( .A(\buff[44][4] ), .B(\buff[45][4] ), .C(\buff[46][4] ), .D(
        \buff[47][4] ), .S0(n9322), .S1(n9325), .Y(n9239) );
  MX4X1 U10840 ( .A(\buff[36][4] ), .B(\buff[37][4] ), .C(\buff[38][4] ), .D(
        \buff[39][4] ), .S0(n9322), .S1(n9325), .Y(n9241) );
  MX4X1 U10841 ( .A(\buff[40][4] ), .B(\buff[41][4] ), .C(\buff[42][4] ), .D(
        \buff[43][4] ), .S0(n9322), .S1(n9328), .Y(n9240) );
  MX4X1 U10842 ( .A(n9262), .B(n9260), .C(n9261), .D(n9259), .S0(n9336), .S1(
        n9334), .Y(n9263) );
  MX4X1 U10843 ( .A(\buff[44][5] ), .B(\buff[45][5] ), .C(\buff[46][5] ), .D(
        \buff[47][5] ), .S0(n9323), .S1(n9328), .Y(n9259) );
  MX4X1 U10844 ( .A(\buff[36][5] ), .B(\buff[37][5] ), .C(\buff[38][5] ), .D(
        \buff[39][5] ), .S0(n9323), .S1(n9328), .Y(n9261) );
  MX4X1 U10845 ( .A(\buff[40][5] ), .B(\buff[41][5] ), .C(\buff[42][5] ), .D(
        \buff[43][5] ), .S0(n9323), .S1(n9328), .Y(n9260) );
  MX4X1 U10846 ( .A(n9282), .B(n9280), .C(n9281), .D(n9279), .S0(n9336), .S1(
        n9334), .Y(n9283) );
  MX4X1 U10847 ( .A(\buff[44][6] ), .B(\buff[45][6] ), .C(\buff[46][6] ), .D(
        \buff[47][6] ), .S0(n9324), .S1(n9329), .Y(n9279) );
  MX4X1 U10848 ( .A(\buff[36][6] ), .B(\buff[37][6] ), .C(\buff[38][6] ), .D(
        \buff[39][6] ), .S0(n9314), .S1(n9330), .Y(n9281) );
  MX4X1 U10849 ( .A(\buff[40][6] ), .B(\buff[41][6] ), .C(\buff[42][6] ), .D(
        \buff[43][6] ), .S0(n9324), .S1(n9329), .Y(n9280) );
  MX4X1 U10850 ( .A(n9302), .B(n9300), .C(n9301), .D(n9299), .S0(n9336), .S1(
        n9333), .Y(n9303) );
  MX4X1 U10851 ( .A(\buff[44][7] ), .B(\buff[45][7] ), .C(\buff[46][7] ), .D(
        \buff[47][7] ), .S0(n9316), .S1(n9331), .Y(n9299) );
  MX4X1 U10852 ( .A(\buff[36][7] ), .B(\buff[37][7] ), .C(\buff[38][7] ), .D(
        \buff[39][7] ), .S0(n9314), .S1(n9331), .Y(n9301) );
  MX4X1 U10853 ( .A(\buff[40][7] ), .B(\buff[41][7] ), .C(\buff[42][7] ), .D(
        \buff[43][7] ), .S0(n9315), .S1(n9331), .Y(n9300) );
  MX4X1 U10854 ( .A(\buff[56][0] ), .B(\buff[57][0] ), .C(\buff[58][0] ), .D(
        \buff[59][0] ), .S0(n9317), .S1(n9329), .Y(n9155) );
  CLKBUFX3 U10855 ( .A(N1657), .Y(n9332) );
  NOR2X1 U10856 ( .A(n9743), .B(n2571), .Y(n2569) );
  CLKBUFX3 U10857 ( .A(N1659), .Y(n9337) );
  CLKBUFX3 U10858 ( .A(N1658), .Y(n9334) );
  NAND2X1 U10859 ( .A(n2574), .B(n2571), .Y(n2563) );
  NAND3X2 U10860 ( .A(n2586), .B(N1656), .C(n2291), .Y(n173) );
  NAND3X2 U10861 ( .A(n2586), .B(N1656), .C(n2132), .Y(n227) );
  NAND3X2 U10862 ( .A(n2586), .B(n2587), .C(n2291), .Y(n186) );
  OAI2BB2XL U10863 ( .B0(n9457), .B1(n138), .A0N(n7291), .A1N(n9457), .Y(n2607) );
  AOI221XL U10864 ( .A0(n9796), .A1(n139), .B0(n9439), .B1(n9430), .C0(n9440), 
        .Y(n138) );
  OAI2BB2XL U10865 ( .B0(n9457), .B1(n142), .A0N(n7321), .A1N(n9457), .Y(n2609) );
  AOI221XL U10866 ( .A0(n9796), .A1(n143), .B0(n9435), .B1(n9430), .C0(n9436), 
        .Y(n142) );
  OAI2BB2XL U10867 ( .B0(n9456), .B1(n156), .A0N(n7315), .A1N(n9456), .Y(n2615) );
  AOI221XL U10868 ( .A0(n9795), .A1(n139), .B0(n9429), .B1(n9439), .C0(n9440), 
        .Y(n156) );
  OAI2BB2XL U10869 ( .B0(n9456), .B1(n157), .A0N(n8356), .A1N(n9456), .Y(n2616) );
  AOI221XL U10870 ( .A0(n9795), .A1(n141), .B0(n9429), .B1(n9437), .C0(n9438), 
        .Y(n157) );
  OAI2BB2XL U10871 ( .B0(n9456), .B1(n158), .A0N(n7249), .A1N(n9456), .Y(n2617) );
  AOI221XL U10872 ( .A0(n9795), .A1(n143), .B0(n9429), .B1(n9435), .C0(n9436), 
        .Y(n158) );
  OAI2BB2XL U10873 ( .B0(n9455), .B1(n170), .A0N(n7339), .A1N(n9455), .Y(n2623) );
  AOI221XL U10874 ( .A0(n9794), .A1(n139), .B0(n9428), .B1(n9439), .C0(n9440), 
        .Y(n170) );
  OAI2BB2XL U10875 ( .B0(n9455), .B1(n171), .A0N(n7388), .A1N(n9455), .Y(n2624) );
  AOI221XL U10876 ( .A0(n9794), .A1(n141), .B0(n9428), .B1(n9437), .C0(n9438), 
        .Y(n171) );
  OAI2BB2XL U10877 ( .B0(n9455), .B1(n172), .A0N(n7391), .A1N(n9455), .Y(n2625) );
  AOI221XL U10878 ( .A0(n9794), .A1(n143), .B0(n9428), .B1(n9435), .C0(n9436), 
        .Y(n172) );
  OAI2BB2XL U10879 ( .B0(n9454), .B1(n183), .A0N(n7364), .A1N(n9454), .Y(n2631) );
  AOI221XL U10880 ( .A0(n9793), .A1(n139), .B0(n9427), .B1(n9439), .C0(n9440), 
        .Y(n183) );
  OAI2BB2XL U10881 ( .B0(n9454), .B1(n184), .A0N(n7294), .A1N(n9454), .Y(n2632) );
  AOI221XL U10882 ( .A0(n9793), .A1(n141), .B0(n9427), .B1(n9437), .C0(n9438), 
        .Y(n184) );
  AOI221XL U10883 ( .A0(n9793), .A1(n143), .B0(n9427), .B1(n9435), .C0(n9436), 
        .Y(n185) );
  OAI2BB2XL U10884 ( .B0(n9453), .B1(n196), .A0N(n7385), .A1N(n9453), .Y(n2639) );
  AOI221XL U10885 ( .A0(n9792), .A1(n139), .B0(n9426), .B1(n9439), .C0(n9440), 
        .Y(n196) );
  OAI2BB2XL U10886 ( .B0(n9453), .B1(n197), .A0N(n7412), .A1N(n9453), .Y(n2640) );
  AOI221XL U10887 ( .A0(n9792), .A1(n141), .B0(n9426), .B1(n9437), .C0(n9438), 
        .Y(n197) );
  OAI2BB2XL U10888 ( .B0(n9453), .B1(n198), .A0N(n7415), .A1N(n9453), .Y(n2641) );
  AOI221XL U10889 ( .A0(n9792), .A1(n143), .B0(n9426), .B1(n9435), .C0(n9436), 
        .Y(n198) );
  OAI2BB2XL U10890 ( .B0(n9452), .B1(n209), .A0N(n7409), .A1N(n9452), .Y(n2647) );
  AOI221XL U10891 ( .A0(n9791), .A1(n139), .B0(n9425), .B1(n9439), .C0(n9440), 
        .Y(n209) );
  OAI2BB2XL U10892 ( .B0(n9452), .B1(n210), .A0N(n7342), .A1N(n9452), .Y(n2648) );
  AOI221XL U10893 ( .A0(n9791), .A1(n141), .B0(n9425), .B1(n9437), .C0(n9438), 
        .Y(n210) );
  OAI2BB2XL U10894 ( .B0(n9452), .B1(n211), .A0N(n7345), .A1N(n9452), .Y(n2649) );
  AOI221XL U10895 ( .A0(n9791), .A1(n143), .B0(n9425), .B1(n9435), .C0(n9436), 
        .Y(n211) );
  OAI2BB2XL U10896 ( .B0(n9451), .B1(n224), .A0N(n7433), .A1N(n9451), .Y(n2655) );
  AOI221XL U10897 ( .A0(n9790), .A1(n139), .B0(n9424), .B1(n9439), .C0(n9440), 
        .Y(n224) );
  OAI2BB2XL U10898 ( .B0(n9451), .B1(n225), .A0N(n7270), .A1N(n9451), .Y(n2656) );
  AOI221XL U10899 ( .A0(n9790), .A1(n141), .B0(n9424), .B1(n9437), .C0(n9438), 
        .Y(n225) );
  OAI2BB2XL U10900 ( .B0(n9451), .B1(n226), .A0N(n7273), .A1N(n9451), .Y(n2657) );
  AOI221XL U10901 ( .A0(n9790), .A1(n143), .B0(n9424), .B1(n9435), .C0(n9436), 
        .Y(n226) );
  OAI221XL U10902 ( .A0(n301), .A1(n302), .B0(n9709), .B1(n9654), .C0(n7455), 
        .Y(n2666) );
  AOI211X1 U10903 ( .A0(n9796), .A1(n9482), .B0(n306), .C0(n307), .Y(n301) );
  OAI222XL U10904 ( .A0(n9429), .A1(n9601), .B0(n311), .B1(n9506), .C0(n9420), 
        .C1(n9597), .Y(n306) );
  OAI221XL U10905 ( .A0(n314), .A1(n302), .B0(n9709), .B1(n9649), .C0(n7457), 
        .Y(n2667) );
  AOI211X1 U10906 ( .A0(n9796), .A1(n9478), .B0(n317), .C0(n318), .Y(n314) );
  OAI222XL U10907 ( .A0(n9429), .A1(n9592), .B0(n311), .B1(n9503), .C0(n9420), 
        .C1(n9588), .Y(n317) );
  OAI221XL U10908 ( .A0(n322), .A1(n302), .B0(n9709), .B1(n9643), .C0(n7459), 
        .Y(n2668) );
  AOI211X1 U10909 ( .A0(n9796), .A1(n9475), .B0(n325), .C0(n326), .Y(n322) );
  OAI222XL U10910 ( .A0(n9429), .A1(n9583), .B0(n311), .B1(n9500), .C0(n9420), 
        .C1(n9579), .Y(n325) );
  OAI221XL U10911 ( .A0(n330), .A1(n302), .B0(n9709), .B1(n9640), .C0(n7461), 
        .Y(n2669) );
  AOI211X1 U10912 ( .A0(n9796), .A1(n9472), .B0(n333), .C0(n334), .Y(n330) );
  OAI222XL U10913 ( .A0(n9429), .A1(n9574), .B0(n311), .B1(n9496), .C0(n9420), 
        .C1(n9570), .Y(n333) );
  OAI221XL U10914 ( .A0(n338), .A1(n302), .B0(n9709), .B1(n9633), .C0(n7463), 
        .Y(n2670) );
  AOI211X1 U10915 ( .A0(n9796), .A1(n9469), .B0(n341), .C0(n342), .Y(n338) );
  OAI222XL U10916 ( .A0(n9429), .A1(n9564), .B0(n311), .B1(n9493), .C0(n9420), 
        .C1(n9562), .Y(n341) );
  OAI221XL U10917 ( .A0(n346), .A1(n302), .B0(n9709), .B1(n9627), .C0(n7465), 
        .Y(n2671) );
  AOI211X1 U10918 ( .A0(n9796), .A1(n9466), .B0(n349), .C0(n350), .Y(n346) );
  OAI222XL U10919 ( .A0(n9429), .A1(n9556), .B0(n311), .B1(n9490), .C0(n9420), 
        .C1(n9552), .Y(n349) );
  AOI211X1 U10920 ( .A0(n9796), .A1(n9463), .B0(n357), .C0(n358), .Y(n354) );
  OAI222XL U10921 ( .A0(n9429), .A1(n9546), .B0(n311), .B1(n9488), .C0(n9420), 
        .C1(n9543), .Y(n357) );
  AOI211X1 U10922 ( .A0(n9796), .A1(n9460), .B0(n370), .C0(n371), .Y(n362) );
  OAI222XL U10923 ( .A0(n9429), .A1(n9537), .B0(n311), .B1(n9485), .C0(n9420), 
        .C1(n9534), .Y(n370) );
  OAI221XL U10924 ( .A0(n376), .A1(n377), .B0(n9703), .B1(n9656), .C0(n7471), 
        .Y(n2674) );
  AOI211X1 U10925 ( .A0(n9795), .A1(n9482), .B0(n380), .C0(n381), .Y(n376) );
  OAI222XL U10926 ( .A0(n9428), .A1(n9600), .B0(n383), .B1(n9507), .C0(n9597), 
        .C1(n9419), .Y(n380) );
  OAI221XL U10927 ( .A0(n385), .A1(n377), .B0(n9703), .B1(n9650), .C0(n7473), 
        .Y(n2675) );
  AOI211X1 U10928 ( .A0(n9795), .A1(n9478), .B0(n387), .C0(n388), .Y(n385) );
  OAI222XL U10929 ( .A0(n9428), .A1(n9592), .B0(n383), .B1(n9504), .C0(n9588), 
        .C1(n9419), .Y(n387) );
  AOI211X1 U10930 ( .A0(n9795), .A1(n9475), .B0(n391), .C0(n392), .Y(n389) );
  OAI222XL U10931 ( .A0(n9428), .A1(n9583), .B0(n383), .B1(n9501), .C0(n9579), 
        .C1(n9419), .Y(n391) );
  AOI211X1 U10932 ( .A0(n9795), .A1(n9472), .B0(n395), .C0(n396), .Y(n393) );
  OAI222XL U10933 ( .A0(n9428), .A1(n9574), .B0(n383), .B1(n9497), .C0(n9570), 
        .C1(n9419), .Y(n395) );
  AOI211X1 U10934 ( .A0(n9795), .A1(n9469), .B0(n399), .C0(n400), .Y(n397) );
  OAI222XL U10935 ( .A0(n9428), .A1(n9564), .B0(n383), .B1(n9495), .C0(n9562), 
        .C1(n9419), .Y(n399) );
  AOI211X1 U10936 ( .A0(n9795), .A1(n9466), .B0(n403), .C0(n404), .Y(n401) );
  OAI222XL U10937 ( .A0(n9428), .A1(n9557), .B0(n383), .B1(n9490), .C0(n9552), 
        .C1(n9419), .Y(n403) );
  AOI211X1 U10938 ( .A0(n9795), .A1(n9463), .B0(n407), .C0(n408), .Y(n405) );
  OAI222XL U10939 ( .A0(n9428), .A1(n9546), .B0(n383), .B1(n9488), .C0(n9543), 
        .C1(n9419), .Y(n407) );
  AOI211X1 U10940 ( .A0(n9795), .A1(n9460), .B0(n413), .C0(n414), .Y(n409) );
  OAI222XL U10941 ( .A0(n9428), .A1(n9537), .B0(n383), .B1(n9485), .C0(n9534), 
        .C1(n9419), .Y(n413) );
  OAI221XL U10942 ( .A0(n416), .A1(n417), .B0(n9696), .B1(n9656), .C0(n7488), 
        .Y(n2682) );
  AOI211X1 U10943 ( .A0(n9794), .A1(n9482), .B0(n420), .C0(n421), .Y(n416) );
  OAI222XL U10944 ( .A0(n9427), .A1(n9600), .B0(n423), .B1(n9507), .C0(n9599), 
        .C1(n9418), .Y(n420) );
  AOI211X1 U10945 ( .A0(n9794), .A1(n9478), .B0(n427), .C0(n428), .Y(n425) );
  OAI222XL U10946 ( .A0(n9427), .A1(n9592), .B0(n423), .B1(n9504), .C0(n9590), 
        .C1(n9418), .Y(n427) );
  AOI211X1 U10947 ( .A0(n9794), .A1(n9475), .B0(n431), .C0(n432), .Y(n429) );
  OAI222XL U10948 ( .A0(n9427), .A1(n9583), .B0(n423), .B1(n9501), .C0(n9581), 
        .C1(n9418), .Y(n431) );
  AOI211X1 U10949 ( .A0(n9794), .A1(n9472), .B0(n435), .C0(n436), .Y(n433) );
  OAI222XL U10950 ( .A0(n9427), .A1(n9574), .B0(n423), .B1(n9498), .C0(n9572), 
        .C1(n9418), .Y(n435) );
  AOI211X1 U10951 ( .A0(n9794), .A1(n9469), .B0(n439), .C0(n440), .Y(n437) );
  OAI222XL U10952 ( .A0(n9427), .A1(n9564), .B0(n423), .B1(n9493), .C0(n9563), 
        .C1(n9418), .Y(n439) );
  AOI211X1 U10953 ( .A0(n9794), .A1(n9466), .B0(n443), .C0(n444), .Y(n441) );
  OAI222XL U10954 ( .A0(n9427), .A1(n9555), .B0(n423), .B1(n9490), .C0(n9554), 
        .C1(n9418), .Y(n443) );
  AOI211X1 U10955 ( .A0(n9794), .A1(n9463), .B0(n447), .C0(n448), .Y(n445) );
  OAI222XL U10956 ( .A0(n9427), .A1(n9546), .B0(n423), .B1(n9487), .C0(n9545), 
        .C1(n9418), .Y(n447) );
  AOI211X1 U10957 ( .A0(n9794), .A1(n9460), .B0(n453), .C0(n454), .Y(n449) );
  OAI222XL U10958 ( .A0(n9427), .A1(n9537), .B0(n423), .B1(n9484), .C0(n9536), 
        .C1(n9418), .Y(n453) );
  AOI211X1 U10959 ( .A0(n9793), .A1(n9482), .B0(n460), .C0(n461), .Y(n456) );
  OAI222XL U10960 ( .A0(n9426), .A1(n9602), .B0(n463), .B1(n9507), .C0(n9599), 
        .C1(n9417), .Y(n460) );
  AOI211X1 U10961 ( .A0(n9793), .A1(n9478), .B0(n467), .C0(n468), .Y(n465) );
  OAI222XL U10962 ( .A0(n9426), .A1(n9592), .B0(n463), .B1(n9504), .C0(n321), 
        .C1(n9417), .Y(n467) );
  AOI211X1 U10963 ( .A0(n9793), .A1(n9475), .B0(n471), .C0(n472), .Y(n469) );
  OAI222XL U10964 ( .A0(n9426), .A1(n9583), .B0(n463), .B1(n9501), .C0(n9581), 
        .C1(n9417), .Y(n471) );
  AOI211X1 U10965 ( .A0(n9793), .A1(n9472), .B0(n475), .C0(n476), .Y(n473) );
  OAI222XL U10966 ( .A0(n9426), .A1(n9574), .B0(n463), .B1(n9498), .C0(n9572), 
        .C1(n9417), .Y(n475) );
  AOI211X1 U10967 ( .A0(n9793), .A1(n9469), .B0(n479), .C0(n480), .Y(n477) );
  OAI222XL U10968 ( .A0(n9426), .A1(n9565), .B0(n463), .B1(n9495), .C0(n9563), 
        .C1(n9417), .Y(n479) );
  AOI211X1 U10969 ( .A0(n9793), .A1(n9466), .B0(n483), .C0(n484), .Y(n481) );
  OAI222XL U10970 ( .A0(n9426), .A1(n352), .B0(n463), .B1(n9492), .C0(n9554), 
        .C1(n9417), .Y(n483) );
  AOI211X1 U10971 ( .A0(n9793), .A1(n9463), .B0(n487), .C0(n488), .Y(n485) );
  OAI222XL U10972 ( .A0(n9426), .A1(n9546), .B0(n463), .B1(n9489), .C0(n9545), 
        .C1(n9417), .Y(n487) );
  AOI211X1 U10973 ( .A0(n9793), .A1(n9460), .B0(n493), .C0(n494), .Y(n489) );
  OAI222XL U10974 ( .A0(n9426), .A1(n9537), .B0(n463), .B1(n9486), .C0(n9536), 
        .C1(n9417), .Y(n493) );
  OAI221XL U10975 ( .A0(n496), .A1(n7521), .B0(n9716), .B1(n9656), .C0(n7516), 
        .Y(n2698) );
  AOI211X1 U10976 ( .A0(n9792), .A1(n9482), .B0(n500), .C0(n501), .Y(n496) );
  OAI222XL U10977 ( .A0(n9425), .A1(n9601), .B0(n503), .B1(n9507), .C0(n9599), 
        .C1(n9416), .Y(n500) );
  AOI211X1 U10978 ( .A0(n9792), .A1(n9478), .B0(n507), .C0(n508), .Y(n505) );
  OAI222XL U10979 ( .A0(n9425), .A1(n9592), .B0(n503), .B1(n9504), .C0(n9590), 
        .C1(n9416), .Y(n507) );
  AOI211X1 U10980 ( .A0(n9792), .A1(n9475), .B0(n511), .C0(n512), .Y(n509) );
  OAI222XL U10981 ( .A0(n9425), .A1(n9583), .B0(n503), .B1(n9501), .C0(n9581), 
        .C1(n9416), .Y(n511) );
  AOI211X1 U10982 ( .A0(n9792), .A1(n9472), .B0(n515), .C0(n516), .Y(n513) );
  OAI222XL U10983 ( .A0(n9425), .A1(n9574), .B0(n503), .B1(n9498), .C0(n9572), 
        .C1(n9416), .Y(n515) );
  AOI211X1 U10984 ( .A0(n9792), .A1(n9469), .B0(n519), .C0(n520), .Y(n517) );
  OAI222XL U10985 ( .A0(n9425), .A1(n9564), .B0(n503), .B1(n9495), .C0(n9563), 
        .C1(n9416), .Y(n519) );
  AOI211X1 U10986 ( .A0(n9792), .A1(n9466), .B0(n523), .C0(n524), .Y(n521) );
  OAI222XL U10987 ( .A0(n9425), .A1(n352), .B0(n503), .B1(n9492), .C0(n9554), 
        .C1(n9416), .Y(n523) );
  AOI211X1 U10988 ( .A0(n9792), .A1(n9463), .B0(n527), .C0(n528), .Y(n525) );
  OAI222XL U10989 ( .A0(n9425), .A1(n9546), .B0(n503), .B1(n9489), .C0(n9545), 
        .C1(n9416), .Y(n527) );
  AOI211X1 U10990 ( .A0(n9792), .A1(n9460), .B0(n533), .C0(n534), .Y(n529) );
  OAI222XL U10991 ( .A0(n9425), .A1(n9537), .B0(n503), .B1(n9486), .C0(n9536), 
        .C1(n9416), .Y(n533) );
  OAI221XL U10992 ( .A0(n536), .A1(n7538), .B0(n9683), .B1(n9654), .C0(n7533), 
        .Y(n2706) );
  AOI211X1 U10993 ( .A0(n9791), .A1(n9482), .B0(n540), .C0(n541), .Y(n536) );
  OAI222XL U10994 ( .A0(n9424), .A1(n9600), .B0(n543), .B1(n9507), .C0(n9599), 
        .C1(n9415), .Y(n540) );
  OAI221XL U10995 ( .A0(n545), .A1(n7538), .B0(n9683), .B1(n9650), .C0(n7535), 
        .Y(n2707) );
  AOI211X1 U10996 ( .A0(n9791), .A1(n9478), .B0(n547), .C0(n548), .Y(n545) );
  OAI222XL U10997 ( .A0(n9424), .A1(n9592), .B0(n543), .B1(n9504), .C0(n9590), 
        .C1(n9415), .Y(n547) );
  OAI221XL U10998 ( .A0(n549), .A1(n7538), .B0(n9683), .B1(n9644), .C0(n7537), 
        .Y(n2708) );
  AOI211X1 U10999 ( .A0(n9791), .A1(n9475), .B0(n551), .C0(n552), .Y(n549) );
  OAI222XL U11000 ( .A0(n9424), .A1(n9583), .B0(n543), .B1(n9501), .C0(n9581), 
        .C1(n9415), .Y(n551) );
  AOI211X1 U11001 ( .A0(n9791), .A1(n9472), .B0(n555), .C0(n556), .Y(n553) );
  OAI222XL U11002 ( .A0(n9424), .A1(n9574), .B0(n543), .B1(n9498), .C0(n9572), 
        .C1(n9415), .Y(n555) );
  AOI211X1 U11003 ( .A0(n9791), .A1(n9469), .B0(n559), .C0(n560), .Y(n557) );
  OAI222XL U11004 ( .A0(n9424), .A1(n9564), .B0(n543), .B1(n9495), .C0(n9563), 
        .C1(n9415), .Y(n559) );
  AOI211X1 U11005 ( .A0(n9791), .A1(n9466), .B0(n563), .C0(n564), .Y(n561) );
  OAI222XL U11006 ( .A0(n9424), .A1(n352), .B0(n543), .B1(n9492), .C0(n9554), 
        .C1(n9415), .Y(n563) );
  AOI211X1 U11007 ( .A0(n9791), .A1(n9463), .B0(n567), .C0(n568), .Y(n565) );
  OAI222XL U11008 ( .A0(n9424), .A1(n9546), .B0(n543), .B1(n9489), .C0(n9545), 
        .C1(n9415), .Y(n567) );
  AOI211X1 U11009 ( .A0(n9791), .A1(n9460), .B0(n573), .C0(n574), .Y(n569) );
  OAI222XL U11010 ( .A0(n9424), .A1(n9537), .B0(n543), .B1(n9486), .C0(n9536), 
        .C1(n9415), .Y(n573) );
  OAI221XL U11011 ( .A0(n576), .A1(n577), .B0(n9676), .B1(n9656), .C0(n7550), 
        .Y(n2714) );
  AOI211X1 U11012 ( .A0(n9790), .A1(n9482), .B0(n580), .C0(n581), .Y(n576) );
  OAI222XL U11013 ( .A0(n9421), .A1(n9601), .B0(n583), .B1(n9507), .C0(n9599), 
        .C1(n9414), .Y(n580) );
  AOI211X1 U11014 ( .A0(n9790), .A1(n9478), .B0(n587), .C0(n588), .Y(n585) );
  OAI222XL U11015 ( .A0(n9421), .A1(n9592), .B0(n583), .B1(n9504), .C0(n321), 
        .C1(n9414), .Y(n587) );
  AOI211X1 U11016 ( .A0(n9790), .A1(n9475), .B0(n591), .C0(n592), .Y(n589) );
  OAI222XL U11017 ( .A0(n9421), .A1(n9583), .B0(n583), .B1(n9501), .C0(n9581), 
        .C1(n9414), .Y(n591) );
  AOI211X1 U11018 ( .A0(n9790), .A1(n9472), .B0(n595), .C0(n596), .Y(n593) );
  OAI222XL U11019 ( .A0(n9421), .A1(n9574), .B0(n583), .B1(n9498), .C0(n9572), 
        .C1(n9414), .Y(n595) );
  AOI211X1 U11020 ( .A0(n9790), .A1(n9469), .B0(n599), .C0(n600), .Y(n597) );
  OAI222XL U11021 ( .A0(n9421), .A1(n9566), .B0(n583), .B1(n9495), .C0(n9563), 
        .C1(n9414), .Y(n599) );
  AOI211X1 U11022 ( .A0(n9790), .A1(n9466), .B0(n603), .C0(n604), .Y(n601) );
  OAI222XL U11023 ( .A0(n9421), .A1(n9556), .B0(n583), .B1(n9492), .C0(n9554), 
        .C1(n9414), .Y(n603) );
  AOI211X1 U11024 ( .A0(n9790), .A1(n9463), .B0(n607), .C0(n608), .Y(n605) );
  OAI222XL U11025 ( .A0(n9421), .A1(n9546), .B0(n583), .B1(n9489), .C0(n9545), 
        .C1(n9414), .Y(n607) );
  AOI211X1 U11026 ( .A0(n9790), .A1(n9460), .B0(n615), .C0(n616), .Y(n609) );
  OAI222XL U11027 ( .A0(n9421), .A1(n9537), .B0(n583), .B1(n9486), .C0(n9536), 
        .C1(n9414), .Y(n615) );
  OAI221XL U11028 ( .A0(n668), .A1(n669), .B0(n9708), .B1(n9656), .C0(n7582), 
        .Y(n2730) );
  AOI211X1 U11029 ( .A0(n9755), .A1(n9482), .B0(n672), .C0(n673), .Y(n668) );
  OAI222XL U11030 ( .A0(n9600), .A1(n9419), .B0(n675), .B1(n9507), .C0(n9599), 
        .C1(n9410), .Y(n672) );
  OAI221XL U11031 ( .A0(n677), .A1(n669), .B0(n9708), .B1(n9648), .C0(n7584), 
        .Y(n2731) );
  AOI211X1 U11032 ( .A0(n9755), .A1(n9478), .B0(n679), .C0(n680), .Y(n677) );
  OAI222XL U11033 ( .A0(n9593), .A1(n9419), .B0(n675), .B1(n9504), .C0(n9589), 
        .C1(n9410), .Y(n679) );
  OAI221XL U11034 ( .A0(n681), .A1(n669), .B0(n9708), .B1(n9642), .C0(n7586), 
        .Y(n2732) );
  AOI211X1 U11035 ( .A0(n9755), .A1(n9475), .B0(n683), .C0(n684), .Y(n681) );
  OAI222XL U11036 ( .A0(n9584), .A1(n9419), .B0(n675), .B1(n9501), .C0(n9581), 
        .C1(n9410), .Y(n683) );
  OAI221XL U11037 ( .A0(n685), .A1(n669), .B0(n9708), .B1(n260), .C0(n7588), 
        .Y(n2733) );
  AOI211X1 U11038 ( .A0(n9755), .A1(n9472), .B0(n687), .C0(n688), .Y(n685) );
  OAI222XL U11039 ( .A0(n9575), .A1(n9419), .B0(n675), .B1(n9498), .C0(n9572), 
        .C1(n9410), .Y(n687) );
  OAI221XL U11040 ( .A0(n689), .A1(n669), .B0(n9708), .B1(n9635), .C0(n7590), 
        .Y(n2734) );
  AOI211X1 U11041 ( .A0(n9755), .A1(n9469), .B0(n691), .C0(n692), .Y(n689) );
  OAI222XL U11042 ( .A0(n9565), .A1(n9419), .B0(n675), .B1(n9495), .C0(n9563), 
        .C1(n9410), .Y(n691) );
  OAI221XL U11043 ( .A0(n693), .A1(n669), .B0(n9708), .B1(n9628), .C0(n7592), 
        .Y(n2735) );
  AOI211X1 U11044 ( .A0(n9755), .A1(n9466), .B0(n695), .C0(n696), .Y(n693) );
  OAI222XL U11045 ( .A0(n9555), .A1(n9419), .B0(n675), .B1(n9492), .C0(n9554), 
        .C1(n9410), .Y(n695) );
  OAI221XL U11046 ( .A0(n697), .A1(n669), .B0(n9708), .B1(n9624), .C0(n7705), 
        .Y(n2736) );
  AOI211X1 U11047 ( .A0(n9755), .A1(n9463), .B0(n699), .C0(n700), .Y(n697) );
  OAI222XL U11048 ( .A0(n9547), .A1(n9419), .B0(n675), .B1(n9489), .C0(n9545), 
        .C1(n9410), .Y(n699) );
  OAI221XL U11049 ( .A0(n701), .A1(n669), .B0(n9708), .B1(n9618), .C0(n7707), 
        .Y(n2737) );
  AOI211X1 U11050 ( .A0(n9755), .A1(n9460), .B0(n706), .C0(n707), .Y(n701) );
  OAI222XL U11051 ( .A0(n9538), .A1(n9419), .B0(n675), .B1(n9486), .C0(n9536), 
        .C1(n9410), .Y(n706) );
  OAI221XL U11052 ( .A0(n709), .A1(n710), .B0(n9702), .B1(n9656), .C0(n7598), 
        .Y(n2738) );
  AOI211X1 U11053 ( .A0(n9754), .A1(n9482), .B0(n713), .C0(n714), .Y(n709) );
  OAI222XL U11054 ( .A0(n9602), .A1(n9418), .B0(n716), .B1(n9507), .C0(n9599), 
        .C1(n9409), .Y(n713) );
  OAI221XL U11055 ( .A0(n718), .A1(n710), .B0(n9702), .B1(n9650), .C0(n7600), 
        .Y(n2739) );
  AOI211X1 U11056 ( .A0(n9754), .A1(n9478), .B0(n720), .C0(n721), .Y(n718) );
  OAI222XL U11057 ( .A0(n9591), .A1(n9418), .B0(n716), .B1(n9504), .C0(n9590), 
        .C1(n9409), .Y(n720) );
  OAI221XL U11058 ( .A0(n722), .A1(n710), .B0(n9702), .B1(n9644), .C0(n7602), 
        .Y(n2740) );
  AOI211X1 U11059 ( .A0(n9754), .A1(n9475), .B0(n724), .C0(n725), .Y(n722) );
  OAI222XL U11060 ( .A0(n9583), .A1(n9418), .B0(n716), .B1(n9501), .C0(n9581), 
        .C1(n9409), .Y(n724) );
  OAI221XL U11061 ( .A0(n726), .A1(n710), .B0(n9702), .B1(n9641), .C0(n7604), 
        .Y(n2741) );
  AOI211X1 U11062 ( .A0(n9754), .A1(n9472), .B0(n728), .C0(n729), .Y(n726) );
  OAI222XL U11063 ( .A0(n9574), .A1(n9418), .B0(n716), .B1(n9498), .C0(n9572), 
        .C1(n9409), .Y(n728) );
  OAI221XL U11064 ( .A0(n730), .A1(n710), .B0(n9702), .B1(n9635), .C0(n7606), 
        .Y(n2742) );
  AOI211X1 U11065 ( .A0(n9754), .A1(n9469), .B0(n732), .C0(n733), .Y(n730) );
  OAI222XL U11066 ( .A0(n9564), .A1(n9418), .B0(n716), .B1(n9495), .C0(n9563), 
        .C1(n9409), .Y(n732) );
  OAI221XL U11067 ( .A0(n734), .A1(n710), .B0(n9702), .B1(n9629), .C0(n7608), 
        .Y(n2743) );
  AOI211X1 U11068 ( .A0(n9754), .A1(n9466), .B0(n736), .C0(n737), .Y(n734) );
  OAI222XL U11069 ( .A0(n9555), .A1(n9418), .B0(n716), .B1(n9492), .C0(n9554), 
        .C1(n9409), .Y(n736) );
  OAI221XL U11070 ( .A0(n738), .A1(n710), .B0(n9702), .B1(n9624), .C0(n7721), 
        .Y(n2744) );
  AOI211X1 U11071 ( .A0(n9754), .A1(n9463), .B0(n740), .C0(n741), .Y(n738) );
  OAI222XL U11072 ( .A0(n9546), .A1(n9418), .B0(n716), .B1(n9489), .C0(n9545), 
        .C1(n9409), .Y(n740) );
  OAI221XL U11073 ( .A0(n742), .A1(n710), .B0(n9702), .B1(n9618), .C0(n7723), 
        .Y(n2745) );
  AOI211X1 U11074 ( .A0(n9754), .A1(n9460), .B0(n745), .C0(n746), .Y(n742) );
  OAI222XL U11075 ( .A0(n9539), .A1(n9418), .B0(n716), .B1(n9486), .C0(n9536), 
        .C1(n9409), .Y(n745) );
  OAI221XL U11076 ( .A0(n748), .A1(n749), .B0(n9695), .B1(n9656), .C0(n7614), 
        .Y(n2746) );
  AOI211X1 U11077 ( .A0(n9753), .A1(n9482), .B0(n752), .C0(n753), .Y(n748) );
  OAI222XL U11078 ( .A0(n9601), .A1(n9417), .B0(n755), .B1(n9507), .C0(n9599), 
        .C1(n9408), .Y(n752) );
  OAI221XL U11079 ( .A0(n757), .A1(n749), .B0(n9695), .B1(n9650), .C0(n7616), 
        .Y(n2747) );
  AOI211X1 U11080 ( .A0(n9753), .A1(n9478), .B0(n759), .C0(n760), .Y(n757) );
  OAI222XL U11081 ( .A0(n9592), .A1(n9417), .B0(n755), .B1(n9504), .C0(n9590), 
        .C1(n9408), .Y(n759) );
  OAI221XL U11082 ( .A0(n761), .A1(n749), .B0(n9695), .B1(n9644), .C0(n7618), 
        .Y(n2748) );
  AOI211X1 U11083 ( .A0(n9753), .A1(n9475), .B0(n763), .C0(n764), .Y(n761) );
  OAI222XL U11084 ( .A0(n9583), .A1(n9417), .B0(n755), .B1(n9501), .C0(n9581), 
        .C1(n9408), .Y(n763) );
  OAI221XL U11085 ( .A0(n765), .A1(n749), .B0(n9695), .B1(n9641), .C0(n7620), 
        .Y(n2749) );
  AOI211X1 U11086 ( .A0(n9753), .A1(n9472), .B0(n767), .C0(n768), .Y(n765) );
  OAI222XL U11087 ( .A0(n9574), .A1(n9417), .B0(n755), .B1(n9498), .C0(n9572), 
        .C1(n9408), .Y(n767) );
  OAI221XL U11088 ( .A0(n769), .A1(n749), .B0(n9695), .B1(n9633), .C0(n7622), 
        .Y(n2750) );
  AOI211X1 U11089 ( .A0(n9753), .A1(n9469), .B0(n771), .C0(n772), .Y(n769) );
  OAI222XL U11090 ( .A0(n9566), .A1(n9417), .B0(n755), .B1(n9495), .C0(n9563), 
        .C1(n9408), .Y(n771) );
  OAI221XL U11091 ( .A0(n773), .A1(n749), .B0(n9695), .B1(n9629), .C0(n7624), 
        .Y(n2751) );
  AOI211X1 U11092 ( .A0(n9753), .A1(n9466), .B0(n775), .C0(n776), .Y(n773) );
  OAI222XL U11093 ( .A0(n9556), .A1(n9417), .B0(n755), .B1(n9492), .C0(n9554), 
        .C1(n9408), .Y(n775) );
  OAI221XL U11094 ( .A0(n777), .A1(n749), .B0(n9695), .B1(n9626), .C0(n7737), 
        .Y(n2752) );
  AOI211X1 U11095 ( .A0(n9753), .A1(n9463), .B0(n779), .C0(n780), .Y(n777) );
  OAI222XL U11096 ( .A0(n9548), .A1(n9417), .B0(n755), .B1(n9489), .C0(n9545), 
        .C1(n9408), .Y(n779) );
  OAI221XL U11097 ( .A0(n781), .A1(n749), .B0(n9695), .B1(n9620), .C0(n7739), 
        .Y(n2753) );
  AOI211X1 U11098 ( .A0(n9753), .A1(n9460), .B0(n784), .C0(n785), .Y(n781) );
  OAI222XL U11099 ( .A0(n9538), .A1(n9417), .B0(n755), .B1(n9486), .C0(n9536), 
        .C1(n9408), .Y(n784) );
  AOI211X1 U11100 ( .A0(n9752), .A1(n9482), .B0(n791), .C0(n792), .Y(n787) );
  OAI222XL U11101 ( .A0(n9600), .A1(n9416), .B0(n794), .B1(n9507), .C0(n9599), 
        .C1(n9407), .Y(n791) );
  AOI211X1 U11102 ( .A0(n9752), .A1(n9478), .B0(n798), .C0(n799), .Y(n796) );
  OAI222XL U11103 ( .A0(n9592), .A1(n9416), .B0(n794), .B1(n9504), .C0(n321), 
        .C1(n9407), .Y(n798) );
  AOI211X1 U11104 ( .A0(n9752), .A1(n9475), .B0(n802), .C0(n803), .Y(n800) );
  OAI222XL U11105 ( .A0(n9584), .A1(n9416), .B0(n794), .B1(n9501), .C0(n9581), 
        .C1(n9407), .Y(n802) );
  AOI211X1 U11106 ( .A0(n9752), .A1(n9472), .B0(n806), .C0(n807), .Y(n804) );
  OAI222XL U11107 ( .A0(n9575), .A1(n9416), .B0(n794), .B1(n9498), .C0(n9572), 
        .C1(n9407), .Y(n806) );
  AOI211X1 U11108 ( .A0(n9752), .A1(n9469), .B0(n810), .C0(n811), .Y(n808) );
  OAI222XL U11109 ( .A0(n9564), .A1(n9416), .B0(n794), .B1(n9495), .C0(n9563), 
        .C1(n9407), .Y(n810) );
  AOI211X1 U11110 ( .A0(n9752), .A1(n9466), .B0(n814), .C0(n815), .Y(n812) );
  OAI222XL U11111 ( .A0(n9557), .A1(n9416), .B0(n794), .B1(n9492), .C0(n9554), 
        .C1(n9407), .Y(n814) );
  AOI211X1 U11112 ( .A0(n9752), .A1(n9463), .B0(n818), .C0(n819), .Y(n816) );
  OAI222XL U11113 ( .A0(n9548), .A1(n9416), .B0(n794), .B1(n9489), .C0(n9545), 
        .C1(n9407), .Y(n818) );
  AOI211X1 U11114 ( .A0(n9752), .A1(n9460), .B0(n823), .C0(n824), .Y(n820) );
  OAI222XL U11115 ( .A0(n9539), .A1(n9416), .B0(n794), .B1(n9486), .C0(n9536), 
        .C1(n9407), .Y(n823) );
  OAI221XL U11116 ( .A0(n826), .A1(n827), .B0(n9715), .B1(n9656), .C0(n7646), 
        .Y(n2762) );
  AOI211X1 U11117 ( .A0(n9751), .A1(n9482), .B0(n830), .C0(n831), .Y(n826) );
  OAI222XL U11118 ( .A0(n9602), .A1(n9415), .B0(n833), .B1(n9507), .C0(n9599), 
        .C1(n9406), .Y(n830) );
  AOI211X1 U11119 ( .A0(n9751), .A1(n9478), .B0(n837), .C0(n838), .Y(n835) );
  OAI222XL U11120 ( .A0(n9591), .A1(n9415), .B0(n833), .B1(n9504), .C0(n9589), 
        .C1(n9406), .Y(n837) );
  AOI211X1 U11121 ( .A0(n9751), .A1(n9475), .B0(n841), .C0(n842), .Y(n839) );
  OAI222XL U11122 ( .A0(n9582), .A1(n9415), .B0(n833), .B1(n9501), .C0(n9581), 
        .C1(n9406), .Y(n841) );
  AOI211X1 U11123 ( .A0(n9751), .A1(n9472), .B0(n845), .C0(n846), .Y(n843) );
  OAI222XL U11124 ( .A0(n9573), .A1(n9415), .B0(n833), .B1(n9498), .C0(n9572), 
        .C1(n9406), .Y(n845) );
  AOI211X1 U11125 ( .A0(n9751), .A1(n9469), .B0(n849), .C0(n850), .Y(n847) );
  OAI222XL U11126 ( .A0(n9564), .A1(n9415), .B0(n833), .B1(n9495), .C0(n9563), 
        .C1(n9406), .Y(n849) );
  AOI211X1 U11127 ( .A0(n9751), .A1(n9466), .B0(n853), .C0(n854), .Y(n851) );
  OAI222XL U11128 ( .A0(n9557), .A1(n9415), .B0(n833), .B1(n9492), .C0(n9554), 
        .C1(n9406), .Y(n853) );
  AOI211X1 U11129 ( .A0(n9751), .A1(n9463), .B0(n857), .C0(n858), .Y(n855) );
  OAI222XL U11130 ( .A0(n9548), .A1(n9415), .B0(n833), .B1(n9489), .C0(n9545), 
        .C1(n9406), .Y(n857) );
  AOI211X1 U11131 ( .A0(n9751), .A1(n9460), .B0(n862), .C0(n863), .Y(n859) );
  OAI222XL U11132 ( .A0(n9539), .A1(n9415), .B0(n833), .B1(n9486), .C0(n9536), 
        .C1(n9406), .Y(n862) );
  OAI221XL U11133 ( .A0(n865), .A1(n866), .B0(n9682), .B1(n9656), .C0(n7662), 
        .Y(n2770) );
  AOI211X1 U11134 ( .A0(n9750), .A1(n9482), .B0(n869), .C0(n870), .Y(n865) );
  OAI222XL U11135 ( .A0(n9602), .A1(n9414), .B0(n872), .B1(n9506), .C0(n9599), 
        .C1(n9405), .Y(n869) );
  OAI221XL U11136 ( .A0(n874), .A1(n866), .B0(n9682), .B1(n9650), .C0(n7664), 
        .Y(n2771) );
  AOI211X1 U11137 ( .A0(n9750), .A1(n9478), .B0(n876), .C0(n877), .Y(n874) );
  OAI222XL U11138 ( .A0(n9592), .A1(n9414), .B0(n872), .B1(n9503), .C0(n9589), 
        .C1(n9405), .Y(n876) );
  OAI221XL U11139 ( .A0(n878), .A1(n866), .B0(n9682), .B1(n9644), .C0(n7666), 
        .Y(n2772) );
  AOI211X1 U11140 ( .A0(n9750), .A1(n9475), .B0(n880), .C0(n881), .Y(n878) );
  OAI222XL U11141 ( .A0(n9583), .A1(n9414), .B0(n872), .B1(n9500), .C0(n9581), 
        .C1(n9405), .Y(n880) );
  OAI221XL U11142 ( .A0(n882), .A1(n866), .B0(n9682), .B1(n9641), .C0(n7668), 
        .Y(n2773) );
  AOI211X1 U11143 ( .A0(n9750), .A1(n9472), .B0(n884), .C0(n885), .Y(n882) );
  OAI222XL U11144 ( .A0(n9574), .A1(n9414), .B0(n872), .B1(n9497), .C0(n9572), 
        .C1(n9405), .Y(n884) );
  OAI221XL U11145 ( .A0(n886), .A1(n866), .B0(n9682), .B1(n9633), .C0(n7670), 
        .Y(n2774) );
  AOI211X1 U11146 ( .A0(n9750), .A1(n9469), .B0(n888), .C0(n889), .Y(n886) );
  OAI222XL U11147 ( .A0(n9564), .A1(n9414), .B0(n872), .B1(n9494), .C0(n9563), 
        .C1(n9405), .Y(n888) );
  OAI221XL U11148 ( .A0(n890), .A1(n866), .B0(n9682), .B1(n9629), .C0(n7672), 
        .Y(n2775) );
  AOI211X1 U11149 ( .A0(n9750), .A1(n9466), .B0(n892), .C0(n893), .Y(n890) );
  OAI222XL U11150 ( .A0(n9557), .A1(n9414), .B0(n872), .B1(n9492), .C0(n9554), 
        .C1(n9405), .Y(n892) );
  OAI221XL U11151 ( .A0(n894), .A1(n866), .B0(n9682), .B1(n9626), .C0(n7785), 
        .Y(n2776) );
  AOI211X1 U11152 ( .A0(n9750), .A1(n9463), .B0(n896), .C0(n897), .Y(n894) );
  OAI222XL U11153 ( .A0(n9548), .A1(n9414), .B0(n872), .B1(n9488), .C0(n9545), 
        .C1(n9405), .Y(n896) );
  OAI221XL U11154 ( .A0(n898), .A1(n866), .B0(n9682), .B1(n9620), .C0(n7787), 
        .Y(n2777) );
  AOI211X1 U11155 ( .A0(n9750), .A1(n9460), .B0(n901), .C0(n902), .Y(n898) );
  OAI222XL U11156 ( .A0(n9539), .A1(n9414), .B0(n872), .B1(n9485), .C0(n9536), 
        .C1(n9405), .Y(n901) );
  OAI221XL U11157 ( .A0(n904), .A1(n905), .B0(n9675), .B1(n9656), .C0(n7678), 
        .Y(n2778) );
  AOI211X1 U11158 ( .A0(n9749), .A1(n9483), .B0(n908), .C0(n909), .Y(n904) );
  OAI222XL U11159 ( .A0(n9602), .A1(n9533), .B0(n911), .B1(n9507), .C0(n9599), 
        .C1(n9404), .Y(n908) );
  OAI221XL U11160 ( .A0(n913), .A1(n905), .B0(n9675), .B1(n9650), .C0(n7680), 
        .Y(n2779) );
  AOI211X1 U11161 ( .A0(n9749), .A1(n9479), .B0(n915), .C0(n916), .Y(n913) );
  OAI222XL U11162 ( .A0(n9592), .A1(n9532), .B0(n911), .B1(n9504), .C0(n9588), 
        .C1(n9404), .Y(n915) );
  OAI221XL U11163 ( .A0(n917), .A1(n905), .B0(n9675), .B1(n9644), .C0(n7682), 
        .Y(n2780) );
  AOI211X1 U11164 ( .A0(n9749), .A1(n9476), .B0(n919), .C0(n920), .Y(n917) );
  OAI222XL U11165 ( .A0(n9583), .A1(n9532), .B0(n911), .B1(n9501), .C0(n9581), 
        .C1(n9404), .Y(n919) );
  OAI221XL U11166 ( .A0(n921), .A1(n905), .B0(n9675), .B1(n9641), .C0(n7684), 
        .Y(n2781) );
  AOI211X1 U11167 ( .A0(n9749), .A1(n9473), .B0(n923), .C0(n924), .Y(n921) );
  OAI222XL U11168 ( .A0(n9574), .A1(n9532), .B0(n911), .B1(n9498), .C0(n9572), 
        .C1(n9404), .Y(n923) );
  OAI221XL U11169 ( .A0(n925), .A1(n905), .B0(n9675), .B1(n9633), .C0(n7686), 
        .Y(n2782) );
  AOI211X1 U11170 ( .A0(n9749), .A1(n9470), .B0(n927), .C0(n928), .Y(n925) );
  OAI222XL U11171 ( .A0(n9565), .A1(n9532), .B0(n911), .B1(n9495), .C0(n9563), 
        .C1(n9404), .Y(n927) );
  OAI221XL U11172 ( .A0(n929), .A1(n905), .B0(n9675), .B1(n9629), .C0(n7688), 
        .Y(n2783) );
  AOI211X1 U11173 ( .A0(n9749), .A1(n9467), .B0(n931), .C0(n932), .Y(n929) );
  OAI222XL U11174 ( .A0(n9557), .A1(n9532), .B0(n911), .B1(n9492), .C0(n9554), 
        .C1(n9404), .Y(n931) );
  OAI221XL U11175 ( .A0(n933), .A1(n905), .B0(n9675), .B1(n9626), .C0(n7801), 
        .Y(n2784) );
  AOI211X1 U11176 ( .A0(n9749), .A1(n9464), .B0(n935), .C0(n936), .Y(n933) );
  OAI222XL U11177 ( .A0(n9548), .A1(n9532), .B0(n911), .B1(n9489), .C0(n9545), 
        .C1(n9404), .Y(n935) );
  OAI221XL U11178 ( .A0(n937), .A1(n905), .B0(n9675), .B1(n9620), .C0(n7803), 
        .Y(n2785) );
  AOI211X1 U11179 ( .A0(n9749), .A1(n9461), .B0(n941), .C0(n942), .Y(n937) );
  OAI222XL U11180 ( .A0(n9539), .A1(n9532), .B0(n911), .B1(n9486), .C0(n9536), 
        .C1(n9404), .Y(n941) );
  OAI221XL U11181 ( .A0(n988), .A1(n989), .B0(n9707), .B1(n9656), .C0(n7710), 
        .Y(n2794) );
  AOI211X1 U11182 ( .A0(n9780), .A1(n9483), .B0(n992), .C0(n993), .Y(n988) );
  OAI222XL U11183 ( .A0(n9602), .A1(n9409), .B0(n995), .B1(n9507), .C0(n9599), 
        .C1(n9400), .Y(n992) );
  OAI221XL U11184 ( .A0(n997), .A1(n989), .B0(n9707), .B1(n9650), .C0(n7712), 
        .Y(n2795) );
  AOI211X1 U11185 ( .A0(n9780), .A1(n9479), .B0(n999), .C0(n1000), .Y(n997) );
  OAI222XL U11186 ( .A0(n9592), .A1(n9409), .B0(n995), .B1(n9504), .C0(n9589), 
        .C1(n9400), .Y(n999) );
  OAI221XL U11187 ( .A0(n1001), .A1(n989), .B0(n9707), .B1(n9644), .C0(n7714), 
        .Y(n2796) );
  AOI211X1 U11188 ( .A0(n9780), .A1(n9476), .B0(n1003), .C0(n1004), .Y(n1001)
         );
  OAI222XL U11189 ( .A0(n9583), .A1(n9409), .B0(n995), .B1(n9501), .C0(n9581), 
        .C1(n9400), .Y(n1003) );
  OAI221XL U11190 ( .A0(n1005), .A1(n989), .B0(n9707), .B1(n9641), .C0(n7716), 
        .Y(n2797) );
  AOI211X1 U11191 ( .A0(n9780), .A1(n9473), .B0(n1007), .C0(n1008), .Y(n1005)
         );
  OAI222XL U11192 ( .A0(n9574), .A1(n9409), .B0(n995), .B1(n9498), .C0(n9572), 
        .C1(n9400), .Y(n1007) );
  OAI221XL U11193 ( .A0(n1009), .A1(n989), .B0(n9707), .B1(n9633), .C0(n7718), 
        .Y(n2798) );
  AOI211X1 U11194 ( .A0(n9780), .A1(n9470), .B0(n1011), .C0(n1012), .Y(n1009)
         );
  OAI222XL U11195 ( .A0(n9564), .A1(n9409), .B0(n995), .B1(n9495), .C0(n9563), 
        .C1(n9400), .Y(n1011) );
  OAI221XL U11196 ( .A0(n1013), .A1(n989), .B0(n9707), .B1(n9629), .C0(n7720), 
        .Y(n2799) );
  AOI211X1 U11197 ( .A0(n9780), .A1(n9467), .B0(n1015), .C0(n1016), .Y(n1013)
         );
  OAI222XL U11198 ( .A0(n9557), .A1(n9409), .B0(n995), .B1(n9492), .C0(n9554), 
        .C1(n9400), .Y(n1015) );
  AOI211X1 U11199 ( .A0(n9780), .A1(n9464), .B0(n1019), .C0(n1020), .Y(n1017)
         );
  OAI222XL U11200 ( .A0(n9548), .A1(n9409), .B0(n995), .B1(n9489), .C0(n9545), 
        .C1(n9400), .Y(n1019) );
  AOI211X1 U11201 ( .A0(n9780), .A1(n9461), .B0(n1026), .C0(n1027), .Y(n1021)
         );
  OAI222XL U11202 ( .A0(n9539), .A1(n9409), .B0(n995), .B1(n9486), .C0(n9536), 
        .C1(n9400), .Y(n1026) );
  OAI221XL U11203 ( .A0(n1029), .A1(n1030), .B0(n9701), .B1(n9656), .C0(n7726), 
        .Y(n2802) );
  AOI211X1 U11204 ( .A0(n9779), .A1(n9483), .B0(n1033), .C0(n1034), .Y(n1029)
         );
  OAI222XL U11205 ( .A0(n9602), .A1(n9408), .B0(n1036), .B1(n9507), .C0(n9599), 
        .C1(n9399), .Y(n1033) );
  OAI221XL U11206 ( .A0(n1038), .A1(n1030), .B0(n9701), .B1(n9650), .C0(n7728), 
        .Y(n2803) );
  AOI211X1 U11207 ( .A0(n9779), .A1(n9479), .B0(n1040), .C0(n1041), .Y(n1038)
         );
  OAI222XL U11208 ( .A0(n9592), .A1(n9408), .B0(n1036), .B1(n9504), .C0(n9588), 
        .C1(n9399), .Y(n1040) );
  OAI221XL U11209 ( .A0(n1042), .A1(n1030), .B0(n9701), .B1(n9644), .C0(n7730), 
        .Y(n2804) );
  AOI211X1 U11210 ( .A0(n9779), .A1(n9476), .B0(n1044), .C0(n1045), .Y(n1042)
         );
  OAI222XL U11211 ( .A0(n9583), .A1(n9408), .B0(n1036), .B1(n9501), .C0(n9581), 
        .C1(n9399), .Y(n1044) );
  OAI221XL U11212 ( .A0(n1046), .A1(n1030), .B0(n9701), .B1(n9641), .C0(n7732), 
        .Y(n2805) );
  AOI211X1 U11213 ( .A0(n9779), .A1(n9473), .B0(n1048), .C0(n1049), .Y(n1046)
         );
  OAI222XL U11214 ( .A0(n9574), .A1(n9408), .B0(n1036), .B1(n9498), .C0(n9572), 
        .C1(n9399), .Y(n1048) );
  OAI221XL U11215 ( .A0(n1050), .A1(n1030), .B0(n9701), .B1(n9633), .C0(n7734), 
        .Y(n2806) );
  AOI211X1 U11216 ( .A0(n9779), .A1(n9470), .B0(n1052), .C0(n1053), .Y(n1050)
         );
  OAI222XL U11217 ( .A0(n9564), .A1(n9408), .B0(n1036), .B1(n9495), .C0(n9563), 
        .C1(n9399), .Y(n1052) );
  OAI221XL U11218 ( .A0(n1054), .A1(n1030), .B0(n9701), .B1(n9629), .C0(n7736), 
        .Y(n2807) );
  AOI211X1 U11219 ( .A0(n9779), .A1(n9467), .B0(n1056), .C0(n1057), .Y(n1054)
         );
  OAI222XL U11220 ( .A0(n9557), .A1(n9408), .B0(n1036), .B1(n9492), .C0(n9554), 
        .C1(n9399), .Y(n1056) );
  AOI211X1 U11221 ( .A0(n9779), .A1(n9464), .B0(n1060), .C0(n1061), .Y(n1058)
         );
  OAI222XL U11222 ( .A0(n9548), .A1(n9408), .B0(n1036), .B1(n9489), .C0(n9545), 
        .C1(n9399), .Y(n1060) );
  AOI211X1 U11223 ( .A0(n9779), .A1(n9461), .B0(n1065), .C0(n1066), .Y(n1062)
         );
  OAI222XL U11224 ( .A0(n9539), .A1(n9408), .B0(n1036), .B1(n9486), .C0(n9536), 
        .C1(n9399), .Y(n1065) );
  OAI221XL U11225 ( .A0(n1068), .A1(n1069), .B0(n9694), .B1(n9656), .C0(n7742), 
        .Y(n2810) );
  AOI211X1 U11226 ( .A0(n9778), .A1(n9483), .B0(n1072), .C0(n1073), .Y(n1068)
         );
  OAI222XL U11227 ( .A0(n9602), .A1(n9407), .B0(n1075), .B1(n9507), .C0(n9598), 
        .C1(n9398), .Y(n1072) );
  OAI221XL U11228 ( .A0(n1077), .A1(n1069), .B0(n9694), .B1(n9650), .C0(n7744), 
        .Y(n2811) );
  AOI211X1 U11229 ( .A0(n9778), .A1(n9479), .B0(n1079), .C0(n1080), .Y(n1077)
         );
  OAI222XL U11230 ( .A0(n9592), .A1(n9407), .B0(n1075), .B1(n9504), .C0(n9589), 
        .C1(n9398), .Y(n1079) );
  OAI221XL U11231 ( .A0(n1081), .A1(n1069), .B0(n9694), .B1(n9644), .C0(n7746), 
        .Y(n2812) );
  AOI211X1 U11232 ( .A0(n9778), .A1(n9476), .B0(n1083), .C0(n1084), .Y(n1081)
         );
  OAI222XL U11233 ( .A0(n9583), .A1(n9407), .B0(n1075), .B1(n9501), .C0(n9580), 
        .C1(n9398), .Y(n1083) );
  OAI221XL U11234 ( .A0(n1085), .A1(n1069), .B0(n9694), .B1(n9641), .C0(n7748), 
        .Y(n2813) );
  AOI211X1 U11235 ( .A0(n9778), .A1(n9473), .B0(n1087), .C0(n1088), .Y(n1085)
         );
  OAI222XL U11236 ( .A0(n9574), .A1(n9407), .B0(n1075), .B1(n9498), .C0(n9571), 
        .C1(n9398), .Y(n1087) );
  OAI221XL U11237 ( .A0(n1089), .A1(n1069), .B0(n9694), .B1(n9635), .C0(n7750), 
        .Y(n2814) );
  AOI211X1 U11238 ( .A0(n9778), .A1(n9470), .B0(n1091), .C0(n1092), .Y(n1089)
         );
  OAI222XL U11239 ( .A0(n344), .A1(n9407), .B0(n1075), .B1(n9495), .C0(n9561), 
        .C1(n9398), .Y(n1091) );
  OAI221XL U11240 ( .A0(n1093), .A1(n1069), .B0(n9694), .B1(n9629), .C0(n7752), 
        .Y(n2815) );
  AOI211X1 U11241 ( .A0(n9778), .A1(n9467), .B0(n1095), .C0(n1096), .Y(n1093)
         );
  OAI222XL U11242 ( .A0(n9557), .A1(n9407), .B0(n1075), .B1(n9492), .C0(n9553), 
        .C1(n9398), .Y(n1095) );
  AOI211X1 U11243 ( .A0(n9778), .A1(n9464), .B0(n1099), .C0(n1100), .Y(n1097)
         );
  OAI222XL U11244 ( .A0(n9548), .A1(n9407), .B0(n1075), .B1(n9489), .C0(n9544), 
        .C1(n9398), .Y(n1099) );
  AOI211X1 U11245 ( .A0(n9778), .A1(n9461), .B0(n1104), .C0(n1105), .Y(n1101)
         );
  OAI222XL U11246 ( .A0(n9539), .A1(n9407), .B0(n1075), .B1(n9486), .C0(n9535), 
        .C1(n9398), .Y(n1104) );
  AOI211X1 U11247 ( .A0(n9777), .A1(n9483), .B0(n1111), .C0(n1112), .Y(n1107)
         );
  OAI222XL U11248 ( .A0(n9602), .A1(n9406), .B0(n1114), .B1(n9506), .C0(n9598), 
        .C1(n9528), .Y(n1111) );
  AOI211X1 U11249 ( .A0(n9777), .A1(n9479), .B0(n1118), .C0(n1119), .Y(n1116)
         );
  OAI222XL U11250 ( .A0(n9591), .A1(n9406), .B0(n1114), .B1(n9503), .C0(n9589), 
        .C1(n9528), .Y(n1118) );
  AOI211X1 U11251 ( .A0(n9777), .A1(n9476), .B0(n1122), .C0(n1123), .Y(n1120)
         );
  OAI222XL U11252 ( .A0(n9582), .A1(n9406), .B0(n1114), .B1(n9500), .C0(n9580), 
        .C1(n9528), .Y(n1122) );
  AOI211X1 U11253 ( .A0(n9777), .A1(n9473), .B0(n1126), .C0(n1127), .Y(n1124)
         );
  OAI222XL U11254 ( .A0(n9573), .A1(n9406), .B0(n1114), .B1(n9497), .C0(n9571), 
        .C1(n9528), .Y(n1126) );
  AOI211X1 U11255 ( .A0(n9777), .A1(n9470), .B0(n1130), .C0(n1131), .Y(n1128)
         );
  OAI222XL U11256 ( .A0(n9564), .A1(n9406), .B0(n1114), .B1(n9494), .C0(n9561), 
        .C1(n9528), .Y(n1130) );
  AOI211X1 U11257 ( .A0(n9777), .A1(n9467), .B0(n1134), .C0(n1135), .Y(n1132)
         );
  OAI222XL U11258 ( .A0(n9557), .A1(n9406), .B0(n1114), .B1(n9490), .C0(n9553), 
        .C1(n9528), .Y(n1134) );
  AOI211X1 U11259 ( .A0(n9777), .A1(n9464), .B0(n1138), .C0(n1139), .Y(n1136)
         );
  OAI222XL U11260 ( .A0(n9548), .A1(n9406), .B0(n1114), .B1(n9488), .C0(n9544), 
        .C1(n9528), .Y(n1138) );
  AOI211X1 U11261 ( .A0(n9777), .A1(n9461), .B0(n1143), .C0(n1144), .Y(n1140)
         );
  OAI222XL U11262 ( .A0(n9539), .A1(n9406), .B0(n1114), .B1(n9485), .C0(n9535), 
        .C1(n9528), .Y(n1143) );
  OAI221XL U11263 ( .A0(n1146), .A1(n1147), .B0(n9714), .B1(n9656), .C0(n7774), 
        .Y(n2826) );
  AOI211X1 U11264 ( .A0(n9776), .A1(n9483), .B0(n1150), .C0(n1151), .Y(n1146)
         );
  OAI222XL U11265 ( .A0(n9602), .A1(n9405), .B0(n1153), .B1(n9506), .C0(n9598), 
        .C1(n9396), .Y(n1150) );
  OAI221XL U11266 ( .A0(n1155), .A1(n1147), .B0(n9714), .B1(n9650), .C0(n7776), 
        .Y(n2827) );
  AOI211X1 U11267 ( .A0(n9776), .A1(n9479), .B0(n1157), .C0(n1158), .Y(n1155)
         );
  OAI222XL U11268 ( .A0(n9592), .A1(n9405), .B0(n1153), .B1(n9503), .C0(n9589), 
        .C1(n9396), .Y(n1157) );
  AOI211X1 U11269 ( .A0(n9776), .A1(n9476), .B0(n1161), .C0(n1162), .Y(n1159)
         );
  OAI222XL U11270 ( .A0(n328), .A1(n9405), .B0(n1153), .B1(n9500), .C0(n9580), 
        .C1(n9396), .Y(n1161) );
  AOI211X1 U11271 ( .A0(n9776), .A1(n9473), .B0(n1165), .C0(n1166), .Y(n1163)
         );
  OAI222XL U11272 ( .A0(n336), .A1(n9405), .B0(n1153), .B1(n9497), .C0(n9571), 
        .C1(n9396), .Y(n1165) );
  AOI211X1 U11273 ( .A0(n9776), .A1(n9470), .B0(n1169), .C0(n1170), .Y(n1167)
         );
  OAI222XL U11274 ( .A0(n9564), .A1(n9405), .B0(n1153), .B1(n9494), .C0(n345), 
        .C1(n9396), .Y(n1169) );
  AOI211X1 U11275 ( .A0(n9776), .A1(n9467), .B0(n1173), .C0(n1174), .Y(n1171)
         );
  OAI222XL U11276 ( .A0(n9557), .A1(n9405), .B0(n1153), .B1(n9490), .C0(n9553), 
        .C1(n9396), .Y(n1173) );
  AOI211X1 U11277 ( .A0(n9776), .A1(n9464), .B0(n1177), .C0(n1178), .Y(n1175)
         );
  OAI222XL U11278 ( .A0(n9548), .A1(n9405), .B0(n1153), .B1(n9488), .C0(n9544), 
        .C1(n9396), .Y(n1177) );
  AOI211X1 U11279 ( .A0(n9776), .A1(n9461), .B0(n1182), .C0(n1183), .Y(n1179)
         );
  OAI222XL U11280 ( .A0(n9539), .A1(n9405), .B0(n1153), .B1(n9485), .C0(n9535), 
        .C1(n9396), .Y(n1182) );
  OAI221XL U11281 ( .A0(n1185), .A1(n1186), .B0(n9681), .B1(n9656), .C0(n7790), 
        .Y(n2834) );
  AOI211X1 U11282 ( .A0(n9775), .A1(n9483), .B0(n1189), .C0(n1190), .Y(n1185)
         );
  OAI222XL U11283 ( .A0(n9602), .A1(n9404), .B0(n1192), .B1(n9506), .C0(n9598), 
        .C1(n9395), .Y(n1189) );
  OAI221XL U11284 ( .A0(n1194), .A1(n1186), .B0(n9681), .B1(n9650), .C0(n7792), 
        .Y(n2835) );
  AOI211X1 U11285 ( .A0(n9775), .A1(n9479), .B0(n1196), .C0(n1197), .Y(n1194)
         );
  OAI222XL U11286 ( .A0(n9591), .A1(n9404), .B0(n1192), .B1(n9503), .C0(n9589), 
        .C1(n9395), .Y(n1196) );
  OAI221XL U11287 ( .A0(n1198), .A1(n1186), .B0(n9681), .B1(n9644), .C0(n7794), 
        .Y(n2836) );
  AOI211X1 U11288 ( .A0(n9775), .A1(n9476), .B0(n1200), .C0(n1201), .Y(n1198)
         );
  OAI222XL U11289 ( .A0(n9583), .A1(n9404), .B0(n1192), .B1(n9500), .C0(n9580), 
        .C1(n9395), .Y(n1200) );
  OAI221XL U11290 ( .A0(n1202), .A1(n1186), .B0(n9681), .B1(n9641), .C0(n7796), 
        .Y(n2837) );
  AOI211X1 U11291 ( .A0(n9775), .A1(n9473), .B0(n1204), .C0(n1205), .Y(n1202)
         );
  OAI222XL U11292 ( .A0(n9574), .A1(n9404), .B0(n1192), .B1(n9497), .C0(n9571), 
        .C1(n9395), .Y(n1204) );
  OAI221XL U11293 ( .A0(n1206), .A1(n1186), .B0(n9681), .B1(n9634), .C0(n7798), 
        .Y(n2838) );
  AOI211X1 U11294 ( .A0(n9775), .A1(n9470), .B0(n1208), .C0(n1209), .Y(n1206)
         );
  OAI222XL U11295 ( .A0(n344), .A1(n9404), .B0(n1192), .B1(n9494), .C0(n9562), 
        .C1(n9395), .Y(n1208) );
  OAI221XL U11296 ( .A0(n1210), .A1(n1186), .B0(n9681), .B1(n9629), .C0(n7800), 
        .Y(n2839) );
  AOI211X1 U11297 ( .A0(n9775), .A1(n9467), .B0(n1212), .C0(n1213), .Y(n1210)
         );
  OAI222XL U11298 ( .A0(n9557), .A1(n9404), .B0(n1192), .B1(n9492), .C0(n9553), 
        .C1(n9395), .Y(n1212) );
  AOI211X1 U11299 ( .A0(n9775), .A1(n9464), .B0(n1216), .C0(n1217), .Y(n1214)
         );
  OAI222XL U11300 ( .A0(n9548), .A1(n9404), .B0(n1192), .B1(n9488), .C0(n9544), 
        .C1(n9395), .Y(n1216) );
  AOI211X1 U11301 ( .A0(n9775), .A1(n9461), .B0(n1221), .C0(n1222), .Y(n1218)
         );
  OAI222XL U11302 ( .A0(n9539), .A1(n9404), .B0(n1192), .B1(n9485), .C0(n9535), 
        .C1(n9395), .Y(n1221) );
  OAI221XL U11303 ( .A0(n1224), .A1(n1225), .B0(n9674), .B1(n9656), .C0(n7806), 
        .Y(n2842) );
  AOI211X1 U11304 ( .A0(n9774), .A1(n9483), .B0(n1228), .C0(n1229), .Y(n1224)
         );
  OAI222XL U11305 ( .A0(n9602), .A1(n9531), .B0(n1231), .B1(n9506), .C0(n9598), 
        .C1(n9394), .Y(n1228) );
  AOI211X1 U11306 ( .A0(n9774), .A1(n9479), .B0(n1235), .C0(n1236), .Y(n1233)
         );
  OAI222XL U11307 ( .A0(n320), .A1(n9530), .B0(n1231), .B1(n9503), .C0(n9589), 
        .C1(n9394), .Y(n1235) );
  AOI211X1 U11308 ( .A0(n9774), .A1(n9476), .B0(n1239), .C0(n1240), .Y(n1237)
         );
  OAI222XL U11309 ( .A0(n9582), .A1(n9530), .B0(n1231), .B1(n9500), .C0(n9580), 
        .C1(n9394), .Y(n1239) );
  AOI211X1 U11310 ( .A0(n9774), .A1(n9473), .B0(n1243), .C0(n1244), .Y(n1241)
         );
  OAI222XL U11311 ( .A0(n9573), .A1(n9530), .B0(n1231), .B1(n9497), .C0(n9571), 
        .C1(n9394), .Y(n1243) );
  AOI211X1 U11312 ( .A0(n9774), .A1(n9470), .B0(n1247), .C0(n1248), .Y(n1245)
         );
  OAI222XL U11313 ( .A0(n9564), .A1(n9530), .B0(n1231), .B1(n9494), .C0(n345), 
        .C1(n9394), .Y(n1247) );
  AOI211X1 U11314 ( .A0(n9774), .A1(n9467), .B0(n1251), .C0(n1252), .Y(n1249)
         );
  OAI222XL U11315 ( .A0(n9557), .A1(n9530), .B0(n1231), .B1(n9492), .C0(n9553), 
        .C1(n9394), .Y(n1251) );
  AOI211X1 U11316 ( .A0(n9774), .A1(n9464), .B0(n1255), .C0(n1256), .Y(n1253)
         );
  OAI222XL U11317 ( .A0(n9548), .A1(n9530), .B0(n1231), .B1(n9488), .C0(n9544), 
        .C1(n9394), .Y(n1255) );
  AOI211X1 U11318 ( .A0(n9774), .A1(n9461), .B0(n1261), .C0(n1262), .Y(n1257)
         );
  OAI222XL U11319 ( .A0(n9539), .A1(n9530), .B0(n1231), .B1(n9485), .C0(n9535), 
        .C1(n9394), .Y(n1261) );
  OAI221XL U11320 ( .A0(n1303), .A1(n1304), .B0(n9706), .B1(n9656), .C0(n7839), 
        .Y(n2858) );
  AOI211X1 U11321 ( .A0(n9761), .A1(n9483), .B0(n1307), .C0(n1308), .Y(n1303)
         );
  OAI222XL U11322 ( .A0(n9602), .A1(n9399), .B0(n1310), .B1(n9506), .C0(n9598), 
        .C1(n9390), .Y(n1307) );
  OAI221XL U11323 ( .A0(n1312), .A1(n1304), .B0(n9706), .B1(n9650), .C0(n7841), 
        .Y(n2859) );
  AOI211X1 U11324 ( .A0(n9761), .A1(n9479), .B0(n1314), .C0(n1315), .Y(n1312)
         );
  OAI222XL U11325 ( .A0(n9591), .A1(n9399), .B0(n1310), .B1(n9503), .C0(n9589), 
        .C1(n9390), .Y(n1314) );
  OAI221XL U11326 ( .A0(n1316), .A1(n1304), .B0(n9706), .B1(n9644), .C0(n7843), 
        .Y(n2860) );
  AOI211X1 U11327 ( .A0(n9761), .A1(n9476), .B0(n1318), .C0(n1319), .Y(n1316)
         );
  OAI222XL U11328 ( .A0(n9582), .A1(n9399), .B0(n1310), .B1(n9500), .C0(n9580), 
        .C1(n9390), .Y(n1318) );
  OAI221XL U11329 ( .A0(n1320), .A1(n1304), .B0(n9706), .B1(n9641), .C0(n7845), 
        .Y(n2861) );
  AOI211X1 U11330 ( .A0(n9761), .A1(n9473), .B0(n1322), .C0(n1323), .Y(n1320)
         );
  OAI222XL U11331 ( .A0(n336), .A1(n9399), .B0(n1310), .B1(n9497), .C0(n9571), 
        .C1(n9390), .Y(n1322) );
  OAI221XL U11332 ( .A0(n1324), .A1(n1304), .B0(n9706), .B1(n9634), .C0(n7847), 
        .Y(n2862) );
  AOI211X1 U11333 ( .A0(n9761), .A1(n9470), .B0(n1326), .C0(n1327), .Y(n1324)
         );
  OAI222XL U11334 ( .A0(n344), .A1(n9399), .B0(n1310), .B1(n9494), .C0(n9561), 
        .C1(n9390), .Y(n1326) );
  OAI221XL U11335 ( .A0(n1328), .A1(n1304), .B0(n9706), .B1(n9629), .C0(n7849), 
        .Y(n2863) );
  AOI211X1 U11336 ( .A0(n9761), .A1(n9467), .B0(n1330), .C0(n1331), .Y(n1328)
         );
  OAI222XL U11337 ( .A0(n9557), .A1(n9399), .B0(n1310), .B1(n9491), .C0(n9553), 
        .C1(n9390), .Y(n1330) );
  OAI221XL U11338 ( .A0(n1332), .A1(n1304), .B0(n9706), .B1(n9626), .C0(n7866), 
        .Y(n2864) );
  AOI211X1 U11339 ( .A0(n9761), .A1(n9464), .B0(n1334), .C0(n1335), .Y(n1332)
         );
  OAI222XL U11340 ( .A0(n9548), .A1(n9399), .B0(n1310), .B1(n9488), .C0(n9544), 
        .C1(n9390), .Y(n1334) );
  OAI221XL U11341 ( .A0(n1336), .A1(n1304), .B0(n9706), .B1(n9620), .C0(n7868), 
        .Y(n2865) );
  AOI211X1 U11342 ( .A0(n9761), .A1(n9461), .B0(n1341), .C0(n1342), .Y(n1336)
         );
  OAI222XL U11343 ( .A0(n9539), .A1(n9399), .B0(n1310), .B1(n9485), .C0(n9535), 
        .C1(n9390), .Y(n1341) );
  OAI221XL U11344 ( .A0(n1344), .A1(n1345), .B0(n9700), .B1(n9655), .C0(n7855), 
        .Y(n2866) );
  AOI211X1 U11345 ( .A0(n9760), .A1(n9483), .B0(n1348), .C0(n1349), .Y(n1344)
         );
  OAI222XL U11346 ( .A0(n9601), .A1(n9398), .B0(n1351), .B1(n9506), .C0(n9598), 
        .C1(n9389), .Y(n1348) );
  OAI221XL U11347 ( .A0(n1353), .A1(n1345), .B0(n9700), .B1(n246), .C0(n7857), 
        .Y(n2867) );
  AOI211X1 U11348 ( .A0(n9760), .A1(n9479), .B0(n1355), .C0(n1356), .Y(n1353)
         );
  OAI222XL U11349 ( .A0(n320), .A1(n9398), .B0(n1351), .B1(n9503), .C0(n9589), 
        .C1(n9389), .Y(n1355) );
  OAI221XL U11350 ( .A0(n1357), .A1(n1345), .B0(n9700), .B1(n253), .C0(n7859), 
        .Y(n2868) );
  AOI211X1 U11351 ( .A0(n9760), .A1(n9476), .B0(n1359), .C0(n1360), .Y(n1357)
         );
  OAI222XL U11352 ( .A0(n328), .A1(n9398), .B0(n1351), .B1(n9500), .C0(n9580), 
        .C1(n9389), .Y(n1359) );
  OAI221XL U11353 ( .A0(n1361), .A1(n1345), .B0(n9700), .B1(n260), .C0(n7861), 
        .Y(n2869) );
  AOI211X1 U11354 ( .A0(n9760), .A1(n9473), .B0(n1363), .C0(n1364), .Y(n1361)
         );
  OAI222XL U11355 ( .A0(n336), .A1(n9398), .B0(n1351), .B1(n9497), .C0(n9571), 
        .C1(n9389), .Y(n1363) );
  OAI221XL U11356 ( .A0(n1365), .A1(n1345), .B0(n9700), .B1(n9634), .C0(n7863), 
        .Y(n2870) );
  AOI211X1 U11357 ( .A0(n9760), .A1(n9470), .B0(n1367), .C0(n1368), .Y(n1365)
         );
  OAI222XL U11358 ( .A0(n9566), .A1(n9398), .B0(n1351), .B1(n9494), .C0(n9561), 
        .C1(n9389), .Y(n1367) );
  OAI221XL U11359 ( .A0(n1369), .A1(n1345), .B0(n9700), .B1(n9628), .C0(n7865), 
        .Y(n2871) );
  AOI211X1 U11360 ( .A0(n9760), .A1(n9467), .B0(n1371), .C0(n1372), .Y(n1369)
         );
  OAI222XL U11361 ( .A0(n9556), .A1(n9398), .B0(n1351), .B1(n9492), .C0(n9553), 
        .C1(n9389), .Y(n1371) );
  OAI221XL U11362 ( .A0(n1373), .A1(n1345), .B0(n9700), .B1(n9624), .C0(n7978), 
        .Y(n2872) );
  AOI211X1 U11363 ( .A0(n9760), .A1(n9464), .B0(n1375), .C0(n1376), .Y(n1373)
         );
  OAI222XL U11364 ( .A0(n9548), .A1(n9398), .B0(n1351), .B1(n9488), .C0(n9544), 
        .C1(n9389), .Y(n1375) );
  OAI221XL U11365 ( .A0(n1377), .A1(n1345), .B0(n9700), .B1(n9619), .C0(n7980), 
        .Y(n2873) );
  AOI211X1 U11366 ( .A0(n9760), .A1(n9461), .B0(n1380), .C0(n1381), .Y(n1377)
         );
  OAI222XL U11367 ( .A0(n9537), .A1(n9398), .B0(n1351), .B1(n9485), .C0(n9535), 
        .C1(n9389), .Y(n1380) );
  OAI221XL U11368 ( .A0(n1383), .A1(n1384), .B0(n9693), .B1(n9655), .C0(n7871), 
        .Y(n2874) );
  AOI211X1 U11369 ( .A0(n9759), .A1(n9483), .B0(n1387), .C0(n1388), .Y(n1383)
         );
  OAI222XL U11370 ( .A0(n9601), .A1(n9529), .B0(n1390), .B1(n9506), .C0(n9598), 
        .C1(n9388), .Y(n1387) );
  OAI221XL U11371 ( .A0(n1392), .A1(n1384), .B0(n9693), .B1(n246), .C0(n7873), 
        .Y(n2875) );
  AOI211X1 U11372 ( .A0(n9759), .A1(n9479), .B0(n1394), .C0(n1395), .Y(n1392)
         );
  OAI222XL U11373 ( .A0(n320), .A1(n9528), .B0(n1390), .B1(n9503), .C0(n9589), 
        .C1(n9388), .Y(n1394) );
  OAI221XL U11374 ( .A0(n1396), .A1(n1384), .B0(n9693), .B1(n253), .C0(n7875), 
        .Y(n2876) );
  AOI211X1 U11375 ( .A0(n9759), .A1(n9476), .B0(n1398), .C0(n1399), .Y(n1396)
         );
  OAI222XL U11376 ( .A0(n328), .A1(n9528), .B0(n1390), .B1(n9500), .C0(n9580), 
        .C1(n9388), .Y(n1398) );
  OAI221XL U11377 ( .A0(n1400), .A1(n1384), .B0(n9693), .B1(n260), .C0(n7877), 
        .Y(n2877) );
  AOI211X1 U11378 ( .A0(n9759), .A1(n9473), .B0(n1402), .C0(n1403), .Y(n1400)
         );
  OAI222XL U11379 ( .A0(n336), .A1(n9528), .B0(n1390), .B1(n9497), .C0(n9571), 
        .C1(n9388), .Y(n1402) );
  OAI221XL U11380 ( .A0(n1404), .A1(n1384), .B0(n9693), .B1(n9634), .C0(n7879), 
        .Y(n2878) );
  AOI211X1 U11381 ( .A0(n9759), .A1(n9470), .B0(n1406), .C0(n1407), .Y(n1404)
         );
  OAI222XL U11382 ( .A0(n9566), .A1(n9528), .B0(n1390), .B1(n9494), .C0(n9561), 
        .C1(n9388), .Y(n1406) );
  OAI221XL U11383 ( .A0(n1408), .A1(n1384), .B0(n9693), .B1(n9628), .C0(n7881), 
        .Y(n2879) );
  AOI211X1 U11384 ( .A0(n9759), .A1(n9467), .B0(n1410), .C0(n1411), .Y(n1408)
         );
  OAI222XL U11385 ( .A0(n9556), .A1(n9528), .B0(n1390), .B1(n9491), .C0(n9553), 
        .C1(n9388), .Y(n1410) );
  OAI221XL U11386 ( .A0(n1412), .A1(n1384), .B0(n9693), .B1(n9624), .C0(n7366), 
        .Y(n2880) );
  AOI211X1 U11387 ( .A0(n9759), .A1(n9464), .B0(n1414), .C0(n1415), .Y(n1412)
         );
  OAI222XL U11388 ( .A0(n9548), .A1(n9528), .B0(n1390), .B1(n9488), .C0(n9544), 
        .C1(n9388), .Y(n1414) );
  OAI221XL U11389 ( .A0(n1416), .A1(n1384), .B0(n9693), .B1(n9619), .C0(n7368), 
        .Y(n2881) );
  AOI211X1 U11390 ( .A0(n9759), .A1(n9461), .B0(n1419), .C0(n1420), .Y(n1416)
         );
  OAI222XL U11391 ( .A0(n9538), .A1(n9528), .B0(n1390), .B1(n9485), .C0(n9535), 
        .C1(n9388), .Y(n1419) );
  OAI221XL U11392 ( .A0(n1463), .A1(n1464), .B0(n9713), .B1(n9655), .C0(n7903), 
        .Y(n2890) );
  AOI211X1 U11393 ( .A0(n9758), .A1(n9483), .B0(n1467), .C0(n1468), .Y(n1463)
         );
  OAI222XL U11394 ( .A0(n9601), .A1(n9395), .B0(n1470), .B1(n9506), .C0(n9598), 
        .C1(n9781), .Y(n1467) );
  AOI211X1 U11395 ( .A0(n9758), .A1(n9479), .B0(n1474), .C0(n1475), .Y(n1472)
         );
  OAI222XL U11396 ( .A0(n9591), .A1(n9395), .B0(n1470), .B1(n9503), .C0(n9589), 
        .C1(n9781), .Y(n1474) );
  AOI211X1 U11397 ( .A0(n9758), .A1(n9476), .B0(n1478), .C0(n1479), .Y(n1476)
         );
  OAI222XL U11398 ( .A0(n9582), .A1(n9395), .B0(n1470), .B1(n9500), .C0(n9580), 
        .C1(n9781), .Y(n1478) );
  AOI211X1 U11399 ( .A0(n9758), .A1(n9473), .B0(n1482), .C0(n1483), .Y(n1480)
         );
  OAI222XL U11400 ( .A0(n9573), .A1(n9395), .B0(n1470), .B1(n9497), .C0(n9571), 
        .C1(n9781), .Y(n1482) );
  AOI211X1 U11401 ( .A0(n9758), .A1(n9470), .B0(n1486), .C0(n1487), .Y(n1484)
         );
  OAI222XL U11402 ( .A0(n9566), .A1(n9395), .B0(n1470), .B1(n9494), .C0(n345), 
        .C1(n9781), .Y(n1486) );
  AOI211X1 U11403 ( .A0(n9758), .A1(n9467), .B0(n1490), .C0(n1491), .Y(n1488)
         );
  OAI222XL U11404 ( .A0(n9556), .A1(n9395), .B0(n1470), .B1(n9491), .C0(n9553), 
        .C1(n9781), .Y(n1490) );
  AOI211X1 U11405 ( .A0(n9758), .A1(n9464), .B0(n1494), .C0(n1495), .Y(n1492)
         );
  OAI222XL U11406 ( .A0(n9547), .A1(n9395), .B0(n1470), .B1(n9488), .C0(n9544), 
        .C1(n9781), .Y(n1494) );
  AOI211X1 U11407 ( .A0(n9758), .A1(n9461), .B0(n1499), .C0(n1500), .Y(n1496)
         );
  OAI222XL U11408 ( .A0(n373), .A1(n9395), .B0(n1470), .B1(n9485), .C0(n9535), 
        .C1(n9781), .Y(n1499) );
  OAI221XL U11409 ( .A0(n1502), .A1(n1503), .B0(n9680), .B1(n9655), .C0(n7919), 
        .Y(n2898) );
  AOI211X1 U11410 ( .A0(n9757), .A1(n9483), .B0(n1506), .C0(n1507), .Y(n1502)
         );
  OAI222XL U11411 ( .A0(n9601), .A1(n9394), .B0(n1509), .B1(n9506), .C0(n9598), 
        .C1(n9385), .Y(n1506) );
  OAI221XL U11412 ( .A0(n1511), .A1(n1503), .B0(n9680), .B1(n246), .C0(n7921), 
        .Y(n2899) );
  AOI211X1 U11413 ( .A0(n9757), .A1(n9479), .B0(n1513), .C0(n1514), .Y(n1511)
         );
  OAI222XL U11414 ( .A0(n320), .A1(n9394), .B0(n1509), .B1(n9503), .C0(n9589), 
        .C1(n9385), .Y(n1513) );
  OAI221XL U11415 ( .A0(n1515), .A1(n1503), .B0(n9680), .B1(n253), .C0(n7923), 
        .Y(n2900) );
  AOI211X1 U11416 ( .A0(n9757), .A1(n9476), .B0(n1517), .C0(n1518), .Y(n1515)
         );
  OAI222XL U11417 ( .A0(n328), .A1(n9394), .B0(n1509), .B1(n9500), .C0(n9580), 
        .C1(n9385), .Y(n1517) );
  OAI221XL U11418 ( .A0(n1519), .A1(n1503), .B0(n9680), .B1(n260), .C0(n7925), 
        .Y(n2901) );
  AOI211X1 U11419 ( .A0(n9757), .A1(n9473), .B0(n1521), .C0(n1522), .Y(n1519)
         );
  OAI222XL U11420 ( .A0(n336), .A1(n9394), .B0(n1509), .B1(n9497), .C0(n9571), 
        .C1(n9385), .Y(n1521) );
  OAI221XL U11421 ( .A0(n1523), .A1(n1503), .B0(n9680), .B1(n9634), .C0(n7927), 
        .Y(n2902) );
  AOI211X1 U11422 ( .A0(n9757), .A1(n9470), .B0(n1525), .C0(n1526), .Y(n1523)
         );
  OAI222XL U11423 ( .A0(n9566), .A1(n9394), .B0(n1509), .B1(n9494), .C0(n9561), 
        .C1(n9385), .Y(n1525) );
  OAI221XL U11424 ( .A0(n1527), .A1(n1503), .B0(n9680), .B1(n9628), .C0(n7929), 
        .Y(n2903) );
  AOI211X1 U11425 ( .A0(n9757), .A1(n9467), .B0(n1529), .C0(n1530), .Y(n1527)
         );
  OAI222XL U11426 ( .A0(n9556), .A1(n9394), .B0(n1509), .B1(n9492), .C0(n9553), 
        .C1(n9385), .Y(n1529) );
  OAI221XL U11427 ( .A0(n1531), .A1(n1503), .B0(n9680), .B1(n9624), .C0(n8042), 
        .Y(n2904) );
  AOI211X1 U11428 ( .A0(n9757), .A1(n9464), .B0(n1533), .C0(n1534), .Y(n1531)
         );
  OAI222XL U11429 ( .A0(n9548), .A1(n9394), .B0(n1509), .B1(n9488), .C0(n9544), 
        .C1(n9385), .Y(n1533) );
  OAI221XL U11430 ( .A0(n1535), .A1(n1503), .B0(n9680), .B1(n9619), .C0(n8044), 
        .Y(n2905) );
  AOI211X1 U11431 ( .A0(n9757), .A1(n9461), .B0(n1538), .C0(n1539), .Y(n1535)
         );
  OAI222XL U11432 ( .A0(n9539), .A1(n9394), .B0(n1509), .B1(n9485), .C0(n9535), 
        .C1(n9385), .Y(n1538) );
  OAI221XL U11433 ( .A0(n1541), .A1(n1542), .B0(n9673), .B1(n9655), .C0(n7935), 
        .Y(n2906) );
  AOI211X1 U11434 ( .A0(n9756), .A1(n9482), .B0(n1545), .C0(n1546), .Y(n1541)
         );
  OAI222XL U11435 ( .A0(n9601), .A1(n9527), .B0(n1548), .B1(n9506), .C0(n9598), 
        .C1(n9384), .Y(n1545) );
  OAI221XL U11436 ( .A0(n1550), .A1(n1542), .B0(n9673), .B1(n246), .C0(n7937), 
        .Y(n2907) );
  AOI211X1 U11437 ( .A0(n9756), .A1(n9480), .B0(n1552), .C0(n1553), .Y(n1550)
         );
  OAI222XL U11438 ( .A0(n320), .A1(n9526), .B0(n1548), .B1(n9503), .C0(n9589), 
        .C1(n9384), .Y(n1552) );
  OAI221XL U11439 ( .A0(n1554), .A1(n1542), .B0(n9673), .B1(n253), .C0(n7939), 
        .Y(n2908) );
  AOI211X1 U11440 ( .A0(n9756), .A1(n9477), .B0(n1556), .C0(n1557), .Y(n1554)
         );
  OAI222XL U11441 ( .A0(n328), .A1(n9526), .B0(n1548), .B1(n9500), .C0(n9580), 
        .C1(n9384), .Y(n1556) );
  OAI221XL U11442 ( .A0(n1558), .A1(n1542), .B0(n9673), .B1(n260), .C0(n7941), 
        .Y(n2909) );
  AOI211X1 U11443 ( .A0(n9756), .A1(n9474), .B0(n1560), .C0(n1561), .Y(n1558)
         );
  OAI222XL U11444 ( .A0(n336), .A1(n9526), .B0(n1548), .B1(n9497), .C0(n9571), 
        .C1(n9384), .Y(n1560) );
  OAI221XL U11445 ( .A0(n1562), .A1(n1542), .B0(n9673), .B1(n9634), .C0(n7943), 
        .Y(n2910) );
  AOI211X1 U11446 ( .A0(n9756), .A1(n9471), .B0(n1564), .C0(n1565), .Y(n1562)
         );
  OAI222XL U11447 ( .A0(n9566), .A1(n9526), .B0(n1548), .B1(n9494), .C0(n9561), 
        .C1(n9384), .Y(n1564) );
  OAI221XL U11448 ( .A0(n1566), .A1(n1542), .B0(n9673), .B1(n9628), .C0(n7945), 
        .Y(n2911) );
  AOI211X1 U11449 ( .A0(n9756), .A1(n9468), .B0(n1568), .C0(n1569), .Y(n1566)
         );
  OAI222XL U11450 ( .A0(n9556), .A1(n9526), .B0(n1548), .B1(n9491), .C0(n9553), 
        .C1(n9384), .Y(n1568) );
  OAI221XL U11451 ( .A0(n1570), .A1(n1542), .B0(n9673), .B1(n9624), .C0(n7834), 
        .Y(n2912) );
  AOI211X1 U11452 ( .A0(n9756), .A1(n9465), .B0(n1572), .C0(n1573), .Y(n1570)
         );
  OAI222XL U11453 ( .A0(n9548), .A1(n9526), .B0(n1548), .B1(n9488), .C0(n9544), 
        .C1(n9384), .Y(n1572) );
  OAI221XL U11454 ( .A0(n1574), .A1(n1542), .B0(n9673), .B1(n9619), .C0(n7836), 
        .Y(n2913) );
  AOI211X1 U11455 ( .A0(n9756), .A1(n9462), .B0(n1578), .C0(n1579), .Y(n1574)
         );
  OAI222XL U11456 ( .A0(n9537), .A1(n9526), .B0(n1548), .B1(n9485), .C0(n9535), 
        .C1(n9384), .Y(n1578) );
  OAI221XL U11457 ( .A0(n1619), .A1(n1620), .B0(n9705), .B1(n9655), .C0(n7967), 
        .Y(n2922) );
  AOI211X1 U11458 ( .A0(n9788), .A1(n9483), .B0(n1623), .C0(n1624), .Y(n1619)
         );
  OAI222XL U11459 ( .A0(n9601), .A1(n9389), .B0(n1626), .B1(n9506), .C0(n9598), 
        .C1(n9522), .Y(n1623) );
  OAI221XL U11460 ( .A0(n1627), .A1(n1620), .B0(n9705), .B1(n246), .C0(n7969), 
        .Y(n2923) );
  AOI211X1 U11461 ( .A0(n9788), .A1(n9480), .B0(n1629), .C0(n1630), .Y(n1627)
         );
  OAI222XL U11462 ( .A0(n9591), .A1(n9389), .B0(n1626), .B1(n9503), .C0(n9589), 
        .C1(n9522), .Y(n1629) );
  OAI221XL U11463 ( .A0(n1631), .A1(n1620), .B0(n9705), .B1(n253), .C0(n7971), 
        .Y(n2924) );
  AOI211X1 U11464 ( .A0(n9788), .A1(n9477), .B0(n1633), .C0(n1634), .Y(n1631)
         );
  OAI222XL U11465 ( .A0(n328), .A1(n9389), .B0(n1626), .B1(n9500), .C0(n9580), 
        .C1(n9522), .Y(n1633) );
  OAI221XL U11466 ( .A0(n1635), .A1(n1620), .B0(n9705), .B1(n260), .C0(n7973), 
        .Y(n2925) );
  AOI211X1 U11467 ( .A0(n9788), .A1(n9474), .B0(n1637), .C0(n1638), .Y(n1635)
         );
  OAI222XL U11468 ( .A0(n9573), .A1(n9389), .B0(n1626), .B1(n9497), .C0(n9571), 
        .C1(n9522), .Y(n1637) );
  OAI221XL U11469 ( .A0(n1639), .A1(n1620), .B0(n9705), .B1(n9634), .C0(n7975), 
        .Y(n2926) );
  AOI211X1 U11470 ( .A0(n9788), .A1(n9471), .B0(n1641), .C0(n1642), .Y(n1639)
         );
  OAI222XL U11471 ( .A0(n9566), .A1(n9389), .B0(n1626), .B1(n9494), .C0(n9562), 
        .C1(n9522), .Y(n1641) );
  OAI221XL U11472 ( .A0(n1643), .A1(n1620), .B0(n9705), .B1(n9628), .C0(n7977), 
        .Y(n2927) );
  AOI211X1 U11473 ( .A0(n9788), .A1(n9468), .B0(n1645), .C0(n1646), .Y(n1643)
         );
  OAI222XL U11474 ( .A0(n9556), .A1(n9389), .B0(n1626), .B1(n9492), .C0(n9553), 
        .C1(n9522), .Y(n1645) );
  OAI221XL U11475 ( .A0(n1647), .A1(n1620), .B0(n9705), .B1(n9624), .C0(n8090), 
        .Y(n2928) );
  AOI211X1 U11476 ( .A0(n9788), .A1(n9465), .B0(n1649), .C0(n1650), .Y(n1647)
         );
  OAI222XL U11477 ( .A0(n9547), .A1(n9389), .B0(n1626), .B1(n9488), .C0(n9544), 
        .C1(n9522), .Y(n1649) );
  OAI221XL U11478 ( .A0(n1651), .A1(n1620), .B0(n9705), .B1(n9619), .C0(n8092), 
        .Y(n2929) );
  AOI211X1 U11479 ( .A0(n9788), .A1(n9462), .B0(n1656), .C0(n1657), .Y(n1651)
         );
  OAI222XL U11480 ( .A0(n9538), .A1(n9389), .B0(n1626), .B1(n9485), .C0(n9535), 
        .C1(n9522), .Y(n1656) );
  OAI221XL U11481 ( .A0(n1659), .A1(n1660), .B0(n9699), .B1(n9655), .C0(n7983), 
        .Y(n2930) );
  AOI211X1 U11482 ( .A0(n9787), .A1(n9481), .B0(n1663), .C0(n1664), .Y(n1659)
         );
  OAI222XL U11483 ( .A0(n9601), .A1(n9388), .B0(n1666), .B1(n9506), .C0(n9598), 
        .C1(n9381), .Y(n1663) );
  OAI221XL U11484 ( .A0(n1668), .A1(n1660), .B0(n9699), .B1(n246), .C0(n7985), 
        .Y(n2931) );
  AOI211X1 U11485 ( .A0(n9787), .A1(n9480), .B0(n1670), .C0(n1671), .Y(n1668)
         );
  OAI222XL U11486 ( .A0(n9591), .A1(n9388), .B0(n1666), .B1(n9503), .C0(n9589), 
        .C1(n9381), .Y(n1670) );
  OAI221XL U11487 ( .A0(n1672), .A1(n1660), .B0(n9699), .B1(n253), .C0(n7987), 
        .Y(n2932) );
  AOI211X1 U11488 ( .A0(n9787), .A1(n9477), .B0(n1674), .C0(n1675), .Y(n1672)
         );
  OAI222XL U11489 ( .A0(n9582), .A1(n9388), .B0(n1666), .B1(n9501), .C0(n9580), 
        .C1(n9381), .Y(n1674) );
  OAI221XL U11490 ( .A0(n1676), .A1(n1660), .B0(n9699), .B1(n9639), .C0(n7989), 
        .Y(n2933) );
  AOI211X1 U11491 ( .A0(n9787), .A1(n9474), .B0(n1678), .C0(n1679), .Y(n1676)
         );
  OAI222XL U11492 ( .A0(n9573), .A1(n9388), .B0(n1666), .B1(n9496), .C0(n9571), 
        .C1(n9381), .Y(n1678) );
  OAI221XL U11493 ( .A0(n1680), .A1(n1660), .B0(n9699), .B1(n9634), .C0(n7991), 
        .Y(n2934) );
  AOI211X1 U11494 ( .A0(n9787), .A1(n9471), .B0(n1682), .C0(n1683), .Y(n1680)
         );
  OAI222XL U11495 ( .A0(n9566), .A1(n9388), .B0(n1666), .B1(n9493), .C0(n9561), 
        .C1(n9381), .Y(n1682) );
  OAI221XL U11496 ( .A0(n1684), .A1(n1660), .B0(n9699), .B1(n9628), .C0(n7993), 
        .Y(n2935) );
  AOI211X1 U11497 ( .A0(n9787), .A1(n9468), .B0(n1686), .C0(n1687), .Y(n1684)
         );
  OAI222XL U11498 ( .A0(n9556), .A1(n9388), .B0(n1666), .B1(n9491), .C0(n9553), 
        .C1(n9381), .Y(n1686) );
  AOI211X1 U11499 ( .A0(n9787), .A1(n9465), .B0(n1690), .C0(n1691), .Y(n1688)
         );
  OAI222XL U11500 ( .A0(n9546), .A1(n9388), .B0(n1666), .B1(n9487), .C0(n9544), 
        .C1(n9381), .Y(n1690) );
  AOI211X1 U11501 ( .A0(n9787), .A1(n9462), .B0(n1695), .C0(n1696), .Y(n1692)
         );
  OAI222XL U11502 ( .A0(n9537), .A1(n9388), .B0(n1666), .B1(n9486), .C0(n9535), 
        .C1(n9381), .Y(n1695) );
  OAI221XL U11503 ( .A0(n1698), .A1(n1699), .B0(n9692), .B1(n9655), .C0(n7999), 
        .Y(n2938) );
  AOI211X1 U11504 ( .A0(n9786), .A1(n9481), .B0(n1702), .C0(n1703), .Y(n1698)
         );
  OAI222XL U11505 ( .A0(n9601), .A1(n9387), .B0(n1705), .B1(n9507), .C0(n9597), 
        .C1(n9380), .Y(n1702) );
  OAI221XL U11506 ( .A0(n1707), .A1(n1699), .B0(n9692), .B1(n9648), .C0(n8001), 
        .Y(n2939) );
  AOI211X1 U11507 ( .A0(n9786), .A1(n9480), .B0(n1709), .C0(n1710), .Y(n1707)
         );
  OAI222XL U11508 ( .A0(n9591), .A1(n9387), .B0(n1705), .B1(n9504), .C0(n9588), 
        .C1(n9380), .Y(n1709) );
  OAI221XL U11509 ( .A0(n1711), .A1(n1699), .B0(n9692), .B1(n9642), .C0(n8003), 
        .Y(n2940) );
  AOI211X1 U11510 ( .A0(n9786), .A1(n9477), .B0(n1713), .C0(n1714), .Y(n1711)
         );
  OAI222XL U11511 ( .A0(n9582), .A1(n9387), .B0(n1705), .B1(n9500), .C0(n9579), 
        .C1(n9380), .Y(n1713) );
  OAI221XL U11512 ( .A0(n1715), .A1(n1699), .B0(n9692), .B1(n9639), .C0(n8005), 
        .Y(n2941) );
  AOI211X1 U11513 ( .A0(n9786), .A1(n9474), .B0(n1717), .C0(n1718), .Y(n1715)
         );
  OAI222XL U11514 ( .A0(n9573), .A1(n9387), .B0(n1705), .B1(n9496), .C0(n9570), 
        .C1(n9380), .Y(n1717) );
  OAI221XL U11515 ( .A0(n1719), .A1(n1699), .B0(n9692), .B1(n9634), .C0(n8007), 
        .Y(n2942) );
  AOI211X1 U11516 ( .A0(n9786), .A1(n9471), .B0(n1721), .C0(n1722), .Y(n1719)
         );
  OAI222XL U11517 ( .A0(n9566), .A1(n9387), .B0(n1705), .B1(n9493), .C0(n9562), 
        .C1(n9380), .Y(n1721) );
  OAI221XL U11518 ( .A0(n1723), .A1(n1699), .B0(n9692), .B1(n9628), .C0(n8009), 
        .Y(n2943) );
  AOI211X1 U11519 ( .A0(n9786), .A1(n9468), .B0(n1725), .C0(n1726), .Y(n1723)
         );
  OAI222XL U11520 ( .A0(n9556), .A1(n9387), .B0(n1705), .B1(n9491), .C0(n9552), 
        .C1(n9380), .Y(n1725) );
  OAI221XL U11521 ( .A0(n1727), .A1(n1699), .B0(n9692), .B1(n9624), .C0(n8123), 
        .Y(n2944) );
  AOI211X1 U11522 ( .A0(n9786), .A1(n9465), .B0(n1729), .C0(n1730), .Y(n1727)
         );
  OAI222XL U11523 ( .A0(n9546), .A1(n9387), .B0(n1705), .B1(n9806), .C0(n9543), 
        .C1(n9380), .Y(n1729) );
  OAI221XL U11524 ( .A0(n1731), .A1(n1699), .B0(n9692), .B1(n9619), .C0(n8125), 
        .Y(n2945) );
  AOI211X1 U11525 ( .A0(n9786), .A1(n9462), .B0(n1734), .C0(n1735), .Y(n1731)
         );
  OAI222XL U11526 ( .A0(n373), .A1(n9387), .B0(n1705), .B1(n9805), .C0(n9534), 
        .C1(n9380), .Y(n1734) );
  AOI211X1 U11527 ( .A0(n9785), .A1(n9733), .B0(n1741), .C0(n1742), .Y(n1737)
         );
  OAI222XL U11528 ( .A0(n9601), .A1(n9781), .B0(n1744), .B1(n9506), .C0(n9597), 
        .C1(n9379), .Y(n1741) );
  AOI211X1 U11529 ( .A0(n9785), .A1(n9480), .B0(n1748), .C0(n1749), .Y(n1746)
         );
  OAI222XL U11530 ( .A0(n9591), .A1(n9781), .B0(n1744), .B1(n9503), .C0(n9588), 
        .C1(n9379), .Y(n1748) );
  AOI211X1 U11531 ( .A0(n9785), .A1(n9477), .B0(n1752), .C0(n1753), .Y(n1750)
         );
  OAI222XL U11532 ( .A0(n9582), .A1(n9781), .B0(n1744), .B1(n9501), .C0(n9579), 
        .C1(n9379), .Y(n1752) );
  AOI211X1 U11533 ( .A0(n9785), .A1(n9474), .B0(n1756), .C0(n1757), .Y(n1754)
         );
  OAI222XL U11534 ( .A0(n9573), .A1(n9781), .B0(n1744), .B1(n9496), .C0(n9570), 
        .C1(n9379), .Y(n1756) );
  AOI211X1 U11535 ( .A0(n9785), .A1(n9471), .B0(n1760), .C0(n1761), .Y(n1758)
         );
  OAI222XL U11536 ( .A0(n9566), .A1(n9781), .B0(n1744), .B1(n9493), .C0(n9562), 
        .C1(n9379), .Y(n1760) );
  AOI211X1 U11537 ( .A0(n9785), .A1(n9468), .B0(n1764), .C0(n1765), .Y(n1762)
         );
  OAI222XL U11538 ( .A0(n9556), .A1(n9781), .B0(n1744), .B1(n9491), .C0(n9552), 
        .C1(n9379), .Y(n1764) );
  AOI211X1 U11539 ( .A0(n9785), .A1(n9465), .B0(n1768), .C0(n1769), .Y(n1766)
         );
  OAI222XL U11540 ( .A0(n9548), .A1(n9781), .B0(n1744), .B1(n9487), .C0(n9543), 
        .C1(n9379), .Y(n1768) );
  AOI211X1 U11541 ( .A0(n9785), .A1(n9462), .B0(n1773), .C0(n1774), .Y(n1770)
         );
  OAI222XL U11542 ( .A0(n9538), .A1(n9781), .B0(n1744), .B1(n9484), .C0(n9534), 
        .C1(n9379), .Y(n1773) );
  OAI221XL U11543 ( .A0(n1776), .A1(n1777), .B0(n9712), .B1(n9655), .C0(n8031), 
        .Y(n2954) );
  AOI211X1 U11544 ( .A0(n9386), .A1(n9733), .B0(n1780), .C0(n1781), .Y(n1776)
         );
  OAI222XL U11545 ( .A0(n9601), .A1(n9385), .B0(n1783), .B1(n9507), .C0(n9597), 
        .C1(n9378), .Y(n1780) );
  AOI211X1 U11546 ( .A0(n9386), .A1(n9480), .B0(n1787), .C0(n1788), .Y(n1785)
         );
  OAI222XL U11547 ( .A0(n9591), .A1(n9385), .B0(n1783), .B1(n9503), .C0(n9588), 
        .C1(n9378), .Y(n1787) );
  AOI211X1 U11548 ( .A0(n9386), .A1(n9477), .B0(n1791), .C0(n1792), .Y(n1789)
         );
  OAI222XL U11549 ( .A0(n9582), .A1(n9385), .B0(n1783), .B1(n9500), .C0(n9579), 
        .C1(n9378), .Y(n1791) );
  AOI211X1 U11550 ( .A0(n9386), .A1(n9474), .B0(n1795), .C0(n1796), .Y(n1793)
         );
  OAI222XL U11551 ( .A0(n9573), .A1(n9385), .B0(n1783), .B1(n9496), .C0(n9570), 
        .C1(n9378), .Y(n1795) );
  AOI211X1 U11552 ( .A0(n9386), .A1(n9471), .B0(n1799), .C0(n1800), .Y(n1797)
         );
  OAI222XL U11553 ( .A0(n9566), .A1(n9385), .B0(n1783), .B1(n9493), .C0(n9562), 
        .C1(n9378), .Y(n1799) );
  AOI211X1 U11554 ( .A0(n9386), .A1(n9468), .B0(n1803), .C0(n1804), .Y(n1801)
         );
  OAI222XL U11555 ( .A0(n9556), .A1(n9385), .B0(n1783), .B1(n9491), .C0(n9552), 
        .C1(n9378), .Y(n1803) );
  AOI211X1 U11556 ( .A0(n9386), .A1(n9465), .B0(n1807), .C0(n1808), .Y(n1805)
         );
  OAI222XL U11557 ( .A0(n9546), .A1(n9385), .B0(n1783), .B1(n9488), .C0(n9543), 
        .C1(n9378), .Y(n1807) );
  AOI211X1 U11558 ( .A0(n9386), .A1(n9462), .B0(n1812), .C0(n1813), .Y(n1809)
         );
  OAI222XL U11559 ( .A0(n373), .A1(n9385), .B0(n1783), .B1(n9484), .C0(n9534), 
        .C1(n9378), .Y(n1812) );
  OAI221XL U11560 ( .A0(n1817), .A1(n1818), .B0(n9679), .B1(n9655), .C0(n8047), 
        .Y(n2962) );
  AOI211X1 U11561 ( .A0(n9784), .A1(n9733), .B0(n1821), .C0(n1822), .Y(n1817)
         );
  OAI222XL U11562 ( .A0(n9600), .A1(n9384), .B0(n1824), .B1(n9506), .C0(n9597), 
        .C1(n9377), .Y(n1821) );
  OAI221XL U11563 ( .A0(n1826), .A1(n1818), .B0(n9679), .B1(n9648), .C0(n8049), 
        .Y(n2963) );
  AOI211X1 U11564 ( .A0(n9784), .A1(n9480), .B0(n1828), .C0(n1829), .Y(n1826)
         );
  OAI222XL U11565 ( .A0(n9593), .A1(n9384), .B0(n1824), .B1(n9503), .C0(n9588), 
        .C1(n9377), .Y(n1828) );
  OAI221XL U11566 ( .A0(n1830), .A1(n1818), .B0(n9679), .B1(n9642), .C0(n8051), 
        .Y(n2964) );
  AOI211X1 U11567 ( .A0(n9784), .A1(n9477), .B0(n1832), .C0(n1833), .Y(n1830)
         );
  OAI222XL U11568 ( .A0(n9584), .A1(n9384), .B0(n1824), .B1(n9500), .C0(n9579), 
        .C1(n9377), .Y(n1832) );
  OAI221XL U11569 ( .A0(n1834), .A1(n1818), .B0(n9679), .B1(n9639), .C0(n8053), 
        .Y(n2965) );
  AOI211X1 U11570 ( .A0(n9784), .A1(n9474), .B0(n1836), .C0(n1837), .Y(n1834)
         );
  OAI222XL U11571 ( .A0(n9575), .A1(n9384), .B0(n1824), .B1(n9497), .C0(n9570), 
        .C1(n9377), .Y(n1836) );
  OAI221XL U11572 ( .A0(n1838), .A1(n1818), .B0(n9679), .B1(n9634), .C0(n8055), 
        .Y(n2966) );
  AOI211X1 U11573 ( .A0(n9784), .A1(n9471), .B0(n1840), .C0(n1841), .Y(n1838)
         );
  OAI222XL U11574 ( .A0(n9565), .A1(n9384), .B0(n1824), .B1(n9494), .C0(n9562), 
        .C1(n9377), .Y(n1840) );
  OAI221XL U11575 ( .A0(n1842), .A1(n1818), .B0(n9679), .B1(n9628), .C0(n8057), 
        .Y(n2967) );
  AOI211X1 U11576 ( .A0(n9784), .A1(n9468), .B0(n1844), .C0(n1845), .Y(n1842)
         );
  OAI222XL U11577 ( .A0(n9555), .A1(n9384), .B0(n1824), .B1(n9491), .C0(n9552), 
        .C1(n9377), .Y(n1844) );
  OAI221XL U11578 ( .A0(n1846), .A1(n1818), .B0(n9679), .B1(n9624), .C0(n8171), 
        .Y(n2968) );
  AOI211X1 U11579 ( .A0(n9784), .A1(n9465), .B0(n1848), .C0(n1849), .Y(n1846)
         );
  OAI222XL U11580 ( .A0(n9547), .A1(n9384), .B0(n1824), .B1(n9488), .C0(n9543), 
        .C1(n9377), .Y(n1848) );
  OAI221XL U11581 ( .A0(n1850), .A1(n1818), .B0(n9679), .B1(n9619), .C0(n8173), 
        .Y(n2969) );
  AOI211X1 U11582 ( .A0(n9784), .A1(n9462), .B0(n1853), .C0(n1854), .Y(n1850)
         );
  OAI222XL U11583 ( .A0(n9538), .A1(n9384), .B0(n1824), .B1(n9485), .C0(n9534), 
        .C1(n9377), .Y(n1853) );
  OAI221XL U11584 ( .A0(n1856), .A1(n1857), .B0(n9672), .B1(n9655), .C0(n8063), 
        .Y(n2970) );
  AOI211X1 U11585 ( .A0(n9783), .A1(n9733), .B0(n1860), .C0(n1861), .Y(n1856)
         );
  OAI222XL U11586 ( .A0(n9600), .A1(n9525), .B0(n1863), .B1(n9506), .C0(n9597), 
        .C1(n9376), .Y(n1860) );
  OAI221XL U11587 ( .A0(n1865), .A1(n1857), .B0(n9672), .B1(n9648), .C0(n8065), 
        .Y(n2971) );
  AOI211X1 U11588 ( .A0(n9783), .A1(n9480), .B0(n1867), .C0(n1868), .Y(n1865)
         );
  OAI222XL U11589 ( .A0(n9593), .A1(n9524), .B0(n1863), .B1(n9503), .C0(n9588), 
        .C1(n9376), .Y(n1867) );
  OAI221XL U11590 ( .A0(n1869), .A1(n1857), .B0(n9672), .B1(n9642), .C0(n8067), 
        .Y(n2972) );
  AOI211X1 U11591 ( .A0(n9783), .A1(n9477), .B0(n1871), .C0(n1872), .Y(n1869)
         );
  OAI222XL U11592 ( .A0(n9584), .A1(n9524), .B0(n1863), .B1(n9501), .C0(n9579), 
        .C1(n9376), .Y(n1871) );
  OAI221XL U11593 ( .A0(n1873), .A1(n1857), .B0(n9672), .B1(n9639), .C0(n8069), 
        .Y(n2973) );
  AOI211X1 U11594 ( .A0(n9783), .A1(n9474), .B0(n1875), .C0(n1876), .Y(n1873)
         );
  OAI222XL U11595 ( .A0(n9575), .A1(n9524), .B0(n1863), .B1(n9496), .C0(n9570), 
        .C1(n9376), .Y(n1875) );
  OAI221XL U11596 ( .A0(n1877), .A1(n1857), .B0(n9672), .B1(n9634), .C0(n8071), 
        .Y(n2974) );
  AOI211X1 U11597 ( .A0(n9783), .A1(n9471), .B0(n1879), .C0(n1880), .Y(n1877)
         );
  OAI222XL U11598 ( .A0(n9565), .A1(n9524), .B0(n1863), .B1(n9493), .C0(n9562), 
        .C1(n9376), .Y(n1879) );
  OAI221XL U11599 ( .A0(n1881), .A1(n1857), .B0(n9672), .B1(n9628), .C0(n8073), 
        .Y(n2975) );
  AOI211X1 U11600 ( .A0(n9783), .A1(n9468), .B0(n1883), .C0(n1884), .Y(n1881)
         );
  OAI222XL U11601 ( .A0(n9555), .A1(n9524), .B0(n1863), .B1(n9491), .C0(n9552), 
        .C1(n9376), .Y(n1883) );
  AOI211X1 U11602 ( .A0(n9783), .A1(n9465), .B0(n1887), .C0(n1888), .Y(n1885)
         );
  OAI222XL U11603 ( .A0(n9547), .A1(n9524), .B0(n1863), .B1(n9487), .C0(n9543), 
        .C1(n9376), .Y(n1887) );
  AOI211X1 U11604 ( .A0(n9783), .A1(n9462), .B0(n1893), .C0(n1894), .Y(n1889)
         );
  OAI222XL U11605 ( .A0(n9538), .A1(n9524), .B0(n1863), .B1(n9486), .C0(n9534), 
        .C1(n9376), .Y(n1893) );
  OAI221XL U11606 ( .A0(n1976), .A1(n1977), .B0(n9698), .B1(n9654), .C0(n8112), 
        .Y(n2994) );
  AOI211X1 U11607 ( .A0(n9767), .A1(n9481), .B0(n1980), .C0(n1981), .Y(n1976)
         );
  OAI222XL U11608 ( .A0(n9600), .A1(n9380), .B0(n1983), .B1(n9506), .C0(n9597), 
        .C1(n9369), .Y(n1980) );
  AOI211X1 U11609 ( .A0(n9767), .A1(n9480), .B0(n1987), .C0(n1988), .Y(n1985)
         );
  OAI222XL U11610 ( .A0(n9593), .A1(n9380), .B0(n1983), .B1(n9504), .C0(n9588), 
        .C1(n9369), .Y(n1987) );
  AOI211X1 U11611 ( .A0(n9767), .A1(n9477), .B0(n1991), .C0(n1992), .Y(n1989)
         );
  OAI222XL U11612 ( .A0(n9584), .A1(n9380), .B0(n1983), .B1(n9501), .C0(n9579), 
        .C1(n9369), .Y(n1991) );
  AOI211X1 U11613 ( .A0(n9767), .A1(n9474), .B0(n1995), .C0(n1996), .Y(n1993)
         );
  OAI222XL U11614 ( .A0(n9575), .A1(n9380), .B0(n1983), .B1(n9496), .C0(n9570), 
        .C1(n9369), .Y(n1995) );
  AOI211X1 U11615 ( .A0(n9767), .A1(n9471), .B0(n1999), .C0(n2000), .Y(n1997)
         );
  OAI222XL U11616 ( .A0(n9565), .A1(n9380), .B0(n1983), .B1(n9493), .C0(n9562), 
        .C1(n9369), .Y(n1999) );
  AOI211X1 U11617 ( .A0(n9767), .A1(n9468), .B0(n2003), .C0(n2004), .Y(n2001)
         );
  OAI222XL U11618 ( .A0(n9555), .A1(n9380), .B0(n1983), .B1(n9491), .C0(n9552), 
        .C1(n9369), .Y(n2003) );
  AOI211X1 U11619 ( .A0(n9767), .A1(n9465), .B0(n2007), .C0(n2008), .Y(n2005)
         );
  OAI222XL U11620 ( .A0(n9547), .A1(n9380), .B0(n1983), .B1(n9489), .C0(n9543), 
        .C1(n9369), .Y(n2007) );
  AOI211X1 U11621 ( .A0(n9767), .A1(n9462), .B0(n2012), .C0(n2013), .Y(n2009)
         );
  OAI222XL U11622 ( .A0(n9538), .A1(n9380), .B0(n1983), .B1(n9484), .C0(n9534), 
        .C1(n9369), .Y(n2012) );
  OAI221XL U11623 ( .A0(n2015), .A1(n2016), .B0(n9691), .B1(n9654), .C0(n8128), 
        .Y(n3002) );
  AOI211X1 U11624 ( .A0(n9766), .A1(n9481), .B0(n2019), .C0(n2020), .Y(n2015)
         );
  OAI222XL U11625 ( .A0(n9600), .A1(n9379), .B0(n2022), .B1(n9507), .C0(n9598), 
        .C1(n9366), .Y(n2019) );
  OAI221XL U11626 ( .A0(n2024), .A1(n2016), .B0(n9691), .B1(n9649), .C0(n8130), 
        .Y(n3003) );
  AOI211X1 U11627 ( .A0(n9766), .A1(n9480), .B0(n2026), .C0(n2027), .Y(n2024)
         );
  OAI222XL U11628 ( .A0(n9593), .A1(n9379), .B0(n2022), .B1(n9504), .C0(n9589), 
        .C1(n9366), .Y(n2026) );
  OAI221XL U11629 ( .A0(n2028), .A1(n2016), .B0(n9691), .B1(n9643), .C0(n8132), 
        .Y(n3004) );
  AOI211X1 U11630 ( .A0(n9766), .A1(n9477), .B0(n2030), .C0(n2031), .Y(n2028)
         );
  OAI222XL U11631 ( .A0(n9584), .A1(n9379), .B0(n2022), .B1(n9500), .C0(n9580), 
        .C1(n9366), .Y(n2030) );
  OAI221XL U11632 ( .A0(n2032), .A1(n2016), .B0(n9691), .B1(n9640), .C0(n8134), 
        .Y(n3005) );
  AOI211X1 U11633 ( .A0(n9766), .A1(n9474), .B0(n2034), .C0(n2035), .Y(n2032)
         );
  OAI222XL U11634 ( .A0(n9575), .A1(n9379), .B0(n2022), .B1(n9496), .C0(n9571), 
        .C1(n9366), .Y(n2034) );
  OAI221XL U11635 ( .A0(n2036), .A1(n2016), .B0(n9691), .B1(n9633), .C0(n8136), 
        .Y(n3006) );
  AOI211X1 U11636 ( .A0(n9766), .A1(n9471), .B0(n2038), .C0(n2039), .Y(n2036)
         );
  OAI222XL U11637 ( .A0(n9565), .A1(n9379), .B0(n2022), .B1(n9493), .C0(n9562), 
        .C1(n9366), .Y(n2038) );
  OAI221XL U11638 ( .A0(n2040), .A1(n2016), .B0(n9691), .B1(n9627), .C0(n8138), 
        .Y(n3007) );
  AOI211X1 U11639 ( .A0(n9766), .A1(n9468), .B0(n2042), .C0(n2043), .Y(n2040)
         );
  OAI222XL U11640 ( .A0(n9555), .A1(n9379), .B0(n2022), .B1(n9491), .C0(n9553), 
        .C1(n9366), .Y(n2042) );
  OAI221XL U11641 ( .A0(n2044), .A1(n2016), .B0(n9691), .B1(n9625), .C0(n8253), 
        .Y(n3008) );
  AOI211X1 U11642 ( .A0(n9766), .A1(n9465), .B0(n2046), .C0(n2047), .Y(n2044)
         );
  OAI222XL U11643 ( .A0(n9547), .A1(n9379), .B0(n2022), .B1(n9489), .C0(n9544), 
        .C1(n9366), .Y(n2046) );
  OAI221XL U11644 ( .A0(n2048), .A1(n2016), .B0(n9691), .B1(n9618), .C0(n8255), 
        .Y(n3009) );
  AOI211X1 U11645 ( .A0(n9766), .A1(n9462), .B0(n2051), .C0(n2052), .Y(n2048)
         );
  OAI222XL U11646 ( .A0(n9538), .A1(n9379), .B0(n2022), .B1(n9805), .C0(n9535), 
        .C1(n9366), .Y(n2051) );
  AOI211X1 U11647 ( .A0(n9765), .A1(n9481), .B0(n2058), .C0(n2059), .Y(n2054)
         );
  OAI222XL U11648 ( .A0(n9600), .A1(n9378), .B0(n2061), .B1(n9507), .C0(n9597), 
        .C1(n9363), .Y(n2058) );
  AOI211X1 U11649 ( .A0(n9765), .A1(n9480), .B0(n2065), .C0(n2066), .Y(n2063)
         );
  OAI222XL U11650 ( .A0(n9593), .A1(n9378), .B0(n2061), .B1(n9504), .C0(n9588), 
        .C1(n9363), .Y(n2065) );
  AOI211X1 U11651 ( .A0(n9765), .A1(n9477), .B0(n2069), .C0(n2070), .Y(n2067)
         );
  OAI222XL U11652 ( .A0(n9584), .A1(n9378), .B0(n2061), .B1(n9500), .C0(n9579), 
        .C1(n9363), .Y(n2069) );
  AOI211X1 U11653 ( .A0(n9765), .A1(n9474), .B0(n2073), .C0(n2074), .Y(n2071)
         );
  OAI222XL U11654 ( .A0(n9575), .A1(n9378), .B0(n2061), .B1(n9496), .C0(n9570), 
        .C1(n9363), .Y(n2073) );
  AOI211X1 U11655 ( .A0(n9765), .A1(n9471), .B0(n2077), .C0(n2078), .Y(n2075)
         );
  OAI222XL U11656 ( .A0(n9565), .A1(n9378), .B0(n2061), .B1(n9493), .C0(n9562), 
        .C1(n9363), .Y(n2077) );
  AOI211X1 U11657 ( .A0(n9765), .A1(n9468), .B0(n2081), .C0(n2082), .Y(n2079)
         );
  OAI222XL U11658 ( .A0(n9555), .A1(n9378), .B0(n2061), .B1(n9491), .C0(n9552), 
        .C1(n9363), .Y(n2081) );
  AOI211X1 U11659 ( .A0(n9765), .A1(n9465), .B0(n2085), .C0(n2086), .Y(n2083)
         );
  OAI222XL U11660 ( .A0(n9547), .A1(n9378), .B0(n2061), .B1(n9487), .C0(n9543), 
        .C1(n9363), .Y(n2085) );
  AOI211X1 U11661 ( .A0(n9765), .A1(n9462), .B0(n2090), .C0(n2091), .Y(n2087)
         );
  OAI222XL U11662 ( .A0(n9538), .A1(n9378), .B0(n2061), .B1(n9485), .C0(n9534), 
        .C1(n9363), .Y(n2090) );
  OAI221XL U11663 ( .A0(n2093), .A1(n2094), .B0(n9711), .B1(n9654), .C0(n8160), 
        .Y(n3018) );
  AOI211X1 U11664 ( .A0(n9764), .A1(n9481), .B0(n2097), .C0(n2098), .Y(n2093)
         );
  OAI222XL U11665 ( .A0(n9600), .A1(n9377), .B0(n2100), .B1(n9505), .C0(n9597), 
        .C1(n9518), .Y(n2097) );
  AOI211X1 U11666 ( .A0(n9764), .A1(n9480), .B0(n2104), .C0(n2105), .Y(n2102)
         );
  OAI222XL U11667 ( .A0(n9593), .A1(n9377), .B0(n2100), .B1(n9502), .C0(n9588), 
        .C1(n9518), .Y(n2104) );
  AOI211X1 U11668 ( .A0(n9764), .A1(n9477), .B0(n2108), .C0(n2109), .Y(n2106)
         );
  OAI222XL U11669 ( .A0(n9584), .A1(n9377), .B0(n2100), .B1(n9499), .C0(n9579), 
        .C1(n9519), .Y(n2108) );
  AOI211X1 U11670 ( .A0(n9764), .A1(n9474), .B0(n2112), .C0(n2113), .Y(n2110)
         );
  OAI222XL U11671 ( .A0(n9575), .A1(n9377), .B0(n2100), .B1(n9496), .C0(n9570), 
        .C1(n9519), .Y(n2112) );
  AOI211X1 U11672 ( .A0(n9764), .A1(n9471), .B0(n2116), .C0(n2117), .Y(n2114)
         );
  OAI222XL U11673 ( .A0(n9565), .A1(n9377), .B0(n2100), .B1(n9495), .C0(n9562), 
        .C1(n9518), .Y(n2116) );
  AOI211X1 U11674 ( .A0(n9764), .A1(n9468), .B0(n2120), .C0(n2121), .Y(n2118)
         );
  OAI222XL U11675 ( .A0(n9555), .A1(n9377), .B0(n2100), .B1(n9490), .C0(n9552), 
        .C1(n9518), .Y(n2120) );
  AOI211X1 U11676 ( .A0(n9764), .A1(n9465), .B0(n2124), .C0(n2125), .Y(n2122)
         );
  OAI222XL U11677 ( .A0(n9547), .A1(n9377), .B0(n2100), .B1(n9487), .C0(n9543), 
        .C1(n9518), .Y(n2124) );
  AOI211X1 U11678 ( .A0(n9764), .A1(n9462), .B0(n2133), .C0(n2134), .Y(n2126)
         );
  OAI222XL U11679 ( .A0(n9538), .A1(n9377), .B0(n2100), .B1(n9484), .C0(n9534), 
        .C1(n9518), .Y(n2133) );
  OAI221XL U11680 ( .A0(n2136), .A1(n2137), .B0(n9678), .B1(n9654), .C0(n8176), 
        .Y(n3026) );
  AOI211X1 U11681 ( .A0(n9763), .A1(n9481), .B0(n2140), .C0(n2141), .Y(n2136)
         );
  OAI222XL U11682 ( .A0(n9600), .A1(n9376), .B0(n2143), .B1(n9506), .C0(n9597), 
        .C1(n9358), .Y(n2140) );
  OAI221XL U11683 ( .A0(n2145), .A1(n2137), .B0(n9678), .B1(n9649), .C0(n8178), 
        .Y(n3027) );
  AOI211X1 U11684 ( .A0(n9763), .A1(n9480), .B0(n2147), .C0(n2148), .Y(n2145)
         );
  OAI222XL U11685 ( .A0(n9593), .A1(n9376), .B0(n2143), .B1(n9503), .C0(n9588), 
        .C1(n9358), .Y(n2147) );
  OAI221XL U11686 ( .A0(n2149), .A1(n2137), .B0(n9678), .B1(n9643), .C0(n8180), 
        .Y(n3028) );
  AOI211X1 U11687 ( .A0(n9763), .A1(n9477), .B0(n2151), .C0(n2152), .Y(n2149)
         );
  OAI222XL U11688 ( .A0(n9584), .A1(n9376), .B0(n2143), .B1(n9501), .C0(n9579), 
        .C1(n9358), .Y(n2151) );
  OAI221XL U11689 ( .A0(n2153), .A1(n2137), .B0(n9678), .B1(n9640), .C0(n8182), 
        .Y(n3029) );
  AOI211X1 U11690 ( .A0(n9763), .A1(n9474), .B0(n2155), .C0(n2156), .Y(n2153)
         );
  OAI222XL U11691 ( .A0(n9575), .A1(n9376), .B0(n2143), .B1(n9496), .C0(n9570), 
        .C1(n9358), .Y(n2155) );
  OAI221XL U11692 ( .A0(n2157), .A1(n2137), .B0(n9678), .B1(n9633), .C0(n8184), 
        .Y(n3030) );
  AOI211X1 U11693 ( .A0(n9763), .A1(n9471), .B0(n2159), .C0(n2160), .Y(n2157)
         );
  OAI222XL U11694 ( .A0(n9565), .A1(n9376), .B0(n2143), .B1(n9493), .C0(n9562), 
        .C1(n9358), .Y(n2159) );
  OAI221XL U11695 ( .A0(n2161), .A1(n2137), .B0(n9678), .B1(n9627), .C0(n8186), 
        .Y(n3031) );
  AOI211X1 U11696 ( .A0(n9763), .A1(n9468), .B0(n2163), .C0(n2164), .Y(n2161)
         );
  OAI222XL U11697 ( .A0(n9555), .A1(n9376), .B0(n2143), .B1(n9491), .C0(n9552), 
        .C1(n9358), .Y(n2163) );
  OAI221XL U11698 ( .A0(n2165), .A1(n2137), .B0(n9678), .B1(n9625), .C0(n8302), 
        .Y(n3032) );
  AOI211X1 U11699 ( .A0(n9763), .A1(n9465), .B0(n2167), .C0(n2168), .Y(n2165)
         );
  OAI222XL U11700 ( .A0(n9547), .A1(n9376), .B0(n2143), .B1(n9488), .C0(n9543), 
        .C1(n9358), .Y(n2167) );
  OAI221XL U11701 ( .A0(n2169), .A1(n2137), .B0(n9678), .B1(n9618), .C0(n8304), 
        .Y(n3033) );
  AOI211X1 U11702 ( .A0(n9763), .A1(n9462), .B0(n2172), .C0(n2173), .Y(n2169)
         );
  OAI222XL U11703 ( .A0(n9538), .A1(n9376), .B0(n2143), .B1(n9486), .C0(n9534), 
        .C1(n9358), .Y(n2172) );
  OAI221XL U11704 ( .A0(n2175), .A1(n2176), .B0(n9671), .B1(n9654), .C0(n8193), 
        .Y(n3034) );
  AOI211X1 U11705 ( .A0(n9762), .A1(n9481), .B0(n2179), .C0(n2180), .Y(n2175)
         );
  OAI222XL U11706 ( .A0(n9600), .A1(n9521), .B0(n2182), .B1(n9507), .C0(n9597), 
        .C1(n9345), .Y(n2179) );
  OAI221XL U11707 ( .A0(n2184), .A1(n2176), .B0(n9671), .B1(n9649), .C0(n8195), 
        .Y(n3035) );
  AOI211X1 U11708 ( .A0(n9762), .A1(n9480), .B0(n2186), .C0(n2187), .Y(n2184)
         );
  OAI222XL U11709 ( .A0(n9593), .A1(n9520), .B0(n2182), .B1(n9504), .C0(n9588), 
        .C1(n9345), .Y(n2186) );
  OAI221XL U11710 ( .A0(n2188), .A1(n2176), .B0(n9671), .B1(n9643), .C0(n8197), 
        .Y(n3036) );
  AOI211X1 U11711 ( .A0(n9762), .A1(n9477), .B0(n2190), .C0(n2191), .Y(n2188)
         );
  OAI222XL U11712 ( .A0(n9584), .A1(n9520), .B0(n2182), .B1(n9500), .C0(n9579), 
        .C1(n2183), .Y(n2190) );
  OAI221XL U11713 ( .A0(n2192), .A1(n2176), .B0(n9671), .B1(n9640), .C0(n8199), 
        .Y(n3037) );
  AOI211X1 U11714 ( .A0(n9762), .A1(n9472), .B0(n2194), .C0(n2195), .Y(n2192)
         );
  OAI222XL U11715 ( .A0(n9575), .A1(n9520), .B0(n2182), .B1(n9496), .C0(n9570), 
        .C1(n9345), .Y(n2194) );
  OAI221XL U11716 ( .A0(n2196), .A1(n2176), .B0(n9671), .B1(n9633), .C0(n8201), 
        .Y(n3038) );
  AOI211X1 U11717 ( .A0(n9762), .A1(n9470), .B0(n2198), .C0(n2199), .Y(n2196)
         );
  OAI222XL U11718 ( .A0(n9565), .A1(n9520), .B0(n2182), .B1(n9493), .C0(n9562), 
        .C1(n2183), .Y(n2198) );
  OAI221XL U11719 ( .A0(n2200), .A1(n2176), .B0(n9671), .B1(n9627), .C0(n8203), 
        .Y(n3039) );
  AOI211X1 U11720 ( .A0(n9762), .A1(n9467), .B0(n2202), .C0(n2203), .Y(n2200)
         );
  OAI222XL U11721 ( .A0(n9555), .A1(n9520), .B0(n2182), .B1(n9491), .C0(n9552), 
        .C1(n9345), .Y(n2202) );
  OAI221XL U11722 ( .A0(n2204), .A1(n2176), .B0(n9671), .B1(n9625), .C0(n8319), 
        .Y(n3040) );
  AOI211X1 U11723 ( .A0(n9762), .A1(n9465), .B0(n2206), .C0(n2207), .Y(n2204)
         );
  OAI222XL U11724 ( .A0(n9547), .A1(n9520), .B0(n2182), .B1(n9806), .C0(n9543), 
        .C1(n2183), .Y(n2206) );
  AOI211X1 U11725 ( .A0(n9762), .A1(n9462), .B0(n2212), .C0(n2213), .Y(n2208)
         );
  OAI222XL U11726 ( .A0(n9538), .A1(n9520), .B0(n2182), .B1(n9805), .C0(n9534), 
        .C1(n9345), .Y(n2212) );
  AOI211X1 U11727 ( .A0(n9773), .A1(n9481), .B0(n2258), .C0(n2259), .Y(n2254)
         );
  OAI222XL U11728 ( .A0(n9599), .A1(n9372), .B0(n2261), .B1(n9506), .C0(n310), 
        .C1(n9369), .Y(n2258) );
  AOI211X1 U11729 ( .A0(n9773), .A1(n9732), .B0(n2264), .C0(n2265), .Y(n2262)
         );
  OAI222XL U11730 ( .A0(n321), .A1(n9372), .B0(n2261), .B1(n9503), .C0(n9592), 
        .C1(n9369), .Y(n2264) );
  AOI211X1 U11731 ( .A0(n9773), .A1(n9731), .B0(n2268), .C0(n2269), .Y(n2266)
         );
  OAI222XL U11732 ( .A0(n9581), .A1(n9372), .B0(n2261), .B1(n9500), .C0(n9583), 
        .C1(n9369), .Y(n2268) );
  AOI211X1 U11733 ( .A0(n9773), .A1(n9474), .B0(n2272), .C0(n2273), .Y(n2270)
         );
  OAI222XL U11734 ( .A0(n9572), .A1(n9372), .B0(n2261), .B1(n9496), .C0(n9574), 
        .C1(n9369), .Y(n2272) );
  AOI211X1 U11735 ( .A0(n9773), .A1(n9729), .B0(n2276), .C0(n2277), .Y(n2274)
         );
  OAI222XL U11736 ( .A0(n9563), .A1(n9372), .B0(n2261), .B1(n9493), .C0(n344), 
        .C1(n9369), .Y(n2276) );
  AOI211X1 U11737 ( .A0(n9773), .A1(n9728), .B0(n2280), .C0(n2281), .Y(n2278)
         );
  OAI222XL U11738 ( .A0(n9554), .A1(n9372), .B0(n2261), .B1(n9491), .C0(n9555), 
        .C1(n9369), .Y(n2280) );
  AOI211X1 U11739 ( .A0(n9773), .A1(n9464), .B0(n2284), .C0(n2285), .Y(n2282)
         );
  OAI222XL U11740 ( .A0(n9545), .A1(n9372), .B0(n2261), .B1(n9489), .C0(n9546), 
        .C1(n9369), .Y(n2284) );
  AOI211X1 U11741 ( .A0(n9773), .A1(n9726), .B0(n2292), .C0(n2293), .Y(n2286)
         );
  OAI222XL U11742 ( .A0(n9536), .A1(n9372), .B0(n2261), .B1(n9486), .C0(n9537), 
        .C1(n9369), .Y(n2292) );
  OAI221XL U11743 ( .A0(n2295), .A1(n8248), .B0(n9697), .B1(n9654), .C0(n8241), 
        .Y(n3058) );
  AOI211X1 U11744 ( .A0(n9772), .A1(n9482), .B0(n2300), .C0(n2301), .Y(n2295)
         );
  OAI222XL U11745 ( .A0(n9599), .A1(n9370), .B0(n2304), .B1(n9506), .C0(n9600), 
        .C1(n9366), .Y(n2300) );
  OAI221XL U11746 ( .A0(n2305), .A1(n8248), .B0(n9697), .B1(n9649), .C0(n8243), 
        .Y(n3059) );
  AOI211X1 U11747 ( .A0(n9772), .A1(n9478), .B0(n2307), .C0(n2308), .Y(n2305)
         );
  OAI222XL U11748 ( .A0(n9590), .A1(n9370), .B0(n2304), .B1(n9503), .C0(n9593), 
        .C1(n9366), .Y(n2307) );
  OAI221XL U11749 ( .A0(n2309), .A1(n8248), .B0(n9697), .B1(n9643), .C0(n8245), 
        .Y(n3060) );
  AOI211X1 U11750 ( .A0(n9772), .A1(n9475), .B0(n2311), .C0(n2312), .Y(n2309)
         );
  OAI222XL U11751 ( .A0(n9580), .A1(n9370), .B0(n2304), .B1(n9501), .C0(n9584), 
        .C1(n9366), .Y(n2311) );
  OAI221XL U11752 ( .A0(n2313), .A1(n8248), .B0(n9697), .B1(n9640), .C0(n8247), 
        .Y(n3061) );
  AOI211X1 U11753 ( .A0(n9772), .A1(n9473), .B0(n2315), .C0(n2316), .Y(n2313)
         );
  OAI222XL U11754 ( .A0(n9571), .A1(n9370), .B0(n2304), .B1(n9496), .C0(n9575), 
        .C1(n9366), .Y(n2315) );
  AOI211X1 U11755 ( .A0(n9772), .A1(n9471), .B0(n2319), .C0(n2320), .Y(n2317)
         );
  OAI222XL U11756 ( .A0(n9561), .A1(n9370), .B0(n2304), .B1(n9493), .C0(n9565), 
        .C1(n9366), .Y(n2319) );
  AOI211X1 U11757 ( .A0(n9772), .A1(n9466), .B0(n2323), .C0(n2324), .Y(n2321)
         );
  OAI222XL U11758 ( .A0(n9552), .A1(n9370), .B0(n2304), .B1(n9491), .C0(n9555), 
        .C1(n9366), .Y(n2323) );
  OAI221XL U11759 ( .A0(n2325), .A1(n8248), .B0(n9697), .B1(n9625), .C0(n7511), 
        .Y(n3064) );
  AOI211X1 U11760 ( .A0(n9772), .A1(n9465), .B0(n2327), .C0(n2328), .Y(n2325)
         );
  OAI222XL U11761 ( .A0(n9544), .A1(n9370), .B0(n2304), .B1(n9806), .C0(n9547), 
        .C1(n9366), .Y(n2327) );
  OAI221XL U11762 ( .A0(n2329), .A1(n8248), .B0(n9697), .B1(n9618), .C0(n7513), 
        .Y(n3065) );
  AOI211X1 U11763 ( .A0(n9772), .A1(n9462), .B0(n2332), .C0(n2333), .Y(n2329)
         );
  OAI222XL U11764 ( .A0(n9534), .A1(n9370), .B0(n2304), .B1(n9805), .C0(n9538), 
        .C1(n9366), .Y(n2332) );
  OAI221XL U11765 ( .A0(n2335), .A1(n2336), .B0(n9690), .B1(n9654), .C0(n8258), 
        .Y(n3066) );
  AOI211X1 U11766 ( .A0(n9771), .A1(n9483), .B0(n2340), .C0(n2341), .Y(n2335)
         );
  OAI222XL U11767 ( .A0(n313), .A1(n9367), .B0(n2344), .B1(n9507), .C0(n310), 
        .C1(n9363), .Y(n2340) );
  OAI221XL U11768 ( .A0(n2345), .A1(n2336), .B0(n9690), .B1(n9649), .C0(n8260), 
        .Y(n3067) );
  AOI211X1 U11769 ( .A0(n9771), .A1(n9478), .B0(n2347), .C0(n2348), .Y(n2345)
         );
  OAI222XL U11770 ( .A0(n9590), .A1(n9367), .B0(n2344), .B1(n9504), .C0(n9592), 
        .C1(n9363), .Y(n2347) );
  OAI221XL U11771 ( .A0(n2349), .A1(n2336), .B0(n9690), .B1(n9643), .C0(n8262), 
        .Y(n3068) );
  AOI211X1 U11772 ( .A0(n9771), .A1(n9475), .B0(n2351), .C0(n2352), .Y(n2349)
         );
  OAI222XL U11773 ( .A0(n9579), .A1(n9367), .B0(n2344), .B1(n9500), .C0(n9583), 
        .C1(n9363), .Y(n2351) );
  AOI211X1 U11774 ( .A0(n9771), .A1(n9472), .B0(n2355), .C0(n2356), .Y(n2353)
         );
  OAI222XL U11775 ( .A0(n9570), .A1(n9367), .B0(n2344), .B1(n9496), .C0(n9574), 
        .C1(n9363), .Y(n2355) );
  AOI211X1 U11776 ( .A0(n9771), .A1(n9470), .B0(n2359), .C0(n2360), .Y(n2357)
         );
  OAI222XL U11777 ( .A0(n9561), .A1(n9367), .B0(n2344), .B1(n9493), .C0(n344), 
        .C1(n9363), .Y(n2359) );
  AOI211X1 U11778 ( .A0(n9771), .A1(n9466), .B0(n2363), .C0(n2364), .Y(n2361)
         );
  OAI222XL U11779 ( .A0(n353), .A1(n9367), .B0(n2344), .B1(n9491), .C0(n352), 
        .C1(n9363), .Y(n2363) );
  OAI221XL U11780 ( .A0(n2365), .A1(n2336), .B0(n9690), .B1(n9625), .C0(n7898), 
        .Y(n3072) );
  AOI211X1 U11781 ( .A0(n9771), .A1(n9464), .B0(n2367), .C0(n2368), .Y(n2365)
         );
  OAI222XL U11782 ( .A0(n9544), .A1(n9367), .B0(n2344), .B1(n9806), .C0(n9546), 
        .C1(n9363), .Y(n2367) );
  OAI221XL U11783 ( .A0(n2369), .A1(n2336), .B0(n9690), .B1(n9618), .C0(n7900), 
        .Y(n3073) );
  AOI211X1 U11784 ( .A0(n9771), .A1(n9460), .B0(n2372), .C0(n2373), .Y(n2369)
         );
  OAI222XL U11785 ( .A0(n374), .A1(n9367), .B0(n2344), .B1(n9485), .C0(n9537), 
        .C1(n9363), .Y(n2372) );
  AOI211X1 U11786 ( .A0(n9770), .A1(n9733), .B0(n2380), .C0(n2381), .Y(n2375)
         );
  OAI222XL U11787 ( .A0(n9597), .A1(n9364), .B0(n2384), .B1(n9505), .C0(n310), 
        .C1(n9518), .Y(n2380) );
  AOI211X1 U11788 ( .A0(n9770), .A1(n9480), .B0(n2387), .C0(n2388), .Y(n2385)
         );
  OAI222XL U11789 ( .A0(n9590), .A1(n9364), .B0(n2384), .B1(n9502), .C0(n9592), 
        .C1(n9518), .Y(n2387) );
  AOI211X1 U11790 ( .A0(n9770), .A1(n9477), .B0(n2391), .C0(n2392), .Y(n2389)
         );
  OAI222XL U11791 ( .A0(n9580), .A1(n9364), .B0(n2384), .B1(n9499), .C0(n9583), 
        .C1(n9518), .Y(n2391) );
  AOI211X1 U11792 ( .A0(n9770), .A1(n9474), .B0(n2395), .C0(n2396), .Y(n2393)
         );
  OAI222XL U11793 ( .A0(n9570), .A1(n9364), .B0(n2384), .B1(n9496), .C0(n9574), 
        .C1(n9518), .Y(n2395) );
  AOI211X1 U11794 ( .A0(n9770), .A1(n9469), .B0(n2399), .C0(n2400), .Y(n2397)
         );
  OAI222XL U11795 ( .A0(n9563), .A1(n9364), .B0(n2384), .B1(n9495), .C0(n9564), 
        .C1(n9518), .Y(n2399) );
  AOI211X1 U11796 ( .A0(n9770), .A1(n9468), .B0(n2403), .C0(n2404), .Y(n2401)
         );
  OAI222XL U11797 ( .A0(n353), .A1(n9364), .B0(n2384), .B1(n9490), .C0(n9556), 
        .C1(n9518), .Y(n2403) );
  AOI211X1 U11798 ( .A0(n9770), .A1(n9465), .B0(n2407), .C0(n2408), .Y(n2405)
         );
  OAI222XL U11799 ( .A0(n9544), .A1(n9364), .B0(n2384), .B1(n9487), .C0(n9546), 
        .C1(n9518), .Y(n2407) );
  AOI211X1 U11800 ( .A0(n9770), .A1(n9461), .B0(n2413), .C0(n2414), .Y(n2409)
         );
  OAI222XL U11801 ( .A0(n374), .A1(n9364), .B0(n2384), .B1(n9484), .C0(n9537), 
        .C1(n9518), .Y(n2413) );
  OAI221XL U11802 ( .A0(n2455), .A1(n2456), .B0(n9677), .B1(n9654), .C0(n8307), 
        .Y(n3090) );
  AOI211X1 U11803 ( .A0(n9769), .A1(n9481), .B0(n2459), .C0(n2460), .Y(n2455)
         );
  OAI222XL U11804 ( .A0(n9597), .A1(n9359), .B0(n2463), .B1(n9505), .C0(n310), 
        .C1(n2183), .Y(n2459) );
  OAI221XL U11805 ( .A0(n2464), .A1(n2456), .B0(n9677), .B1(n9649), .C0(n8309), 
        .Y(n3091) );
  AOI211X1 U11806 ( .A0(n9769), .A1(n9479), .B0(n2466), .C0(n2467), .Y(n2464)
         );
  OAI222XL U11807 ( .A0(n9590), .A1(n9359), .B0(n2463), .B1(n9502), .C0(n9592), 
        .C1(n9345), .Y(n2466) );
  OAI221XL U11808 ( .A0(n2468), .A1(n2456), .B0(n9677), .B1(n9643), .C0(n8311), 
        .Y(n3092) );
  AOI211X1 U11809 ( .A0(n9769), .A1(n9476), .B0(n2470), .C0(n2471), .Y(n2468)
         );
  OAI222XL U11810 ( .A0(n9580), .A1(n9359), .B0(n2463), .B1(n9499), .C0(n9583), 
        .C1(n2183), .Y(n2470) );
  AOI211X1 U11811 ( .A0(n9769), .A1(n9473), .B0(n2474), .C0(n2475), .Y(n2472)
         );
  OAI222XL U11812 ( .A0(n9571), .A1(n9359), .B0(n2463), .B1(n9498), .C0(n9574), 
        .C1(n9345), .Y(n2474) );
  AOI211X1 U11813 ( .A0(n9769), .A1(n9469), .B0(n2478), .C0(n2479), .Y(n2476)
         );
  OAI222XL U11814 ( .A0(n9561), .A1(n9359), .B0(n2463), .B1(n9494), .C0(n344), 
        .C1(n2183), .Y(n2478) );
  AOI211X1 U11815 ( .A0(n9769), .A1(n9467), .B0(n2482), .C0(n2483), .Y(n2480)
         );
  OAI222XL U11816 ( .A0(n9552), .A1(n9359), .B0(n2463), .B1(n9490), .C0(n9557), 
        .C1(n9345), .Y(n2482) );
  OAI221XL U11817 ( .A0(n2484), .A1(n2456), .B0(n9677), .B1(n9625), .C0(n7466), 
        .Y(n3096) );
  AOI211X1 U11818 ( .A0(n9769), .A1(n9464), .B0(n2486), .C0(n2487), .Y(n2484)
         );
  OAI222XL U11819 ( .A0(n9544), .A1(n9359), .B0(n2463), .B1(n9487), .C0(n9546), 
        .C1(n2183), .Y(n2486) );
  OAI221XL U11820 ( .A0(n2488), .A1(n2456), .B0(n9677), .B1(n9618), .C0(n7468), 
        .Y(n3097) );
  AOI211X1 U11821 ( .A0(n9769), .A1(n9461), .B0(n2491), .C0(n2492), .Y(n2488)
         );
  OAI222XL U11822 ( .A0(n9534), .A1(n9359), .B0(n2463), .B1(n9484), .C0(n9537), 
        .C1(n9345), .Y(n2491) );
  OAI221XL U11823 ( .A0(n2494), .A1(n2495), .B0(n9670), .B1(n9655), .C0(n8324), 
        .Y(n3098) );
  AOI211X1 U11824 ( .A0(n9768), .A1(n9481), .B0(n2499), .C0(n2500), .Y(n2494)
         );
  OAI222XL U11825 ( .A0(n9601), .A1(n7236), .B0(n9605), .B1(n2503), .C0(n2504), 
        .C1(n9505), .Y(n2499) );
  OAI221XL U11826 ( .A0(n2505), .A1(n2495), .B0(n9670), .B1(n9648), .C0(n8326), 
        .Y(n3099) );
  AOI211X1 U11827 ( .A0(n9768), .A1(n9479), .B0(n2507), .C0(n2508), .Y(n2505)
         );
  OAI222XL U11828 ( .A0(n9591), .A1(n7236), .B0(n9594), .B1(n2503), .C0(n2504), 
        .C1(n9502), .Y(n2507) );
  OAI221XL U11829 ( .A0(n2509), .A1(n2495), .B0(n9670), .B1(n9642), .C0(n8328), 
        .Y(n3100) );
  AOI211X1 U11830 ( .A0(n9768), .A1(n9476), .B0(n2511), .C0(n2512), .Y(n2509)
         );
  OAI222XL U11831 ( .A0(n9582), .A1(n7236), .B0(n9585), .B1(n2503), .C0(n2504), 
        .C1(n9499), .Y(n2511) );
  AOI211X1 U11832 ( .A0(n9768), .A1(n9730), .B0(n2515), .C0(n2516), .Y(n2513)
         );
  OAI222XL U11833 ( .A0(n9573), .A1(n7236), .B0(n9576), .B1(n2503), .C0(n2504), 
        .C1(n9498), .Y(n2515) );
  AOI211X1 U11834 ( .A0(n9768), .A1(n9471), .B0(n2519), .C0(n2520), .Y(n2517)
         );
  OAI222XL U11835 ( .A0(n9566), .A1(n7236), .B0(n9567), .B1(n2503), .C0(n2504), 
        .C1(n9493), .Y(n2519) );
  AOI211X1 U11836 ( .A0(n9768), .A1(n9468), .B0(n2523), .C0(n2524), .Y(n2521)
         );
  OAI222XL U11837 ( .A0(n9556), .A1(n7236), .B0(n9559), .B1(n2503), .C0(n2504), 
        .C1(n9490), .Y(n2523) );
  OAI221XL U11838 ( .A0(n2525), .A1(n2495), .B0(n9670), .B1(n9624), .C0(n7450), 
        .Y(n3104) );
  AOI211X1 U11839 ( .A0(n9768), .A1(n9463), .B0(n2527), .C0(n2528), .Y(n2525)
         );
  OAI222XL U11840 ( .A0(n9547), .A1(n7236), .B0(n9551), .B1(n2503), .C0(n2504), 
        .C1(n9487), .Y(n2527) );
  OAI221XL U11841 ( .A0(n2529), .A1(n2495), .B0(n9670), .B1(n9619), .C0(n7452), 
        .Y(n3105) );
  AOI211X1 U11842 ( .A0(n9768), .A1(n9460), .B0(n2532), .C0(n2533), .Y(n2529)
         );
  OAI222XL U11843 ( .A0(n373), .A1(n7236), .B0(n9541), .B1(n2503), .C0(n2504), 
        .C1(n9484), .Y(n2532) );
  MXI2X1 U11844 ( .A(\buff[25][0] ), .B(\buff[29][0] ), .S0(n8947), .Y(n8644)
         );
  MXI2X1 U11845 ( .A(\buff[25][1] ), .B(\buff[29][1] ), .S0(n8431), .Y(n8657)
         );
  MXI2X1 U11846 ( .A(n8479), .B(n8478), .S0(n8922), .Y(n8740) );
  MX4X1 U11847 ( .A(\buff[8][0] ), .B(\buff[12][0] ), .C(\buff[10][0] ), .D(
        \buff[14][0] ), .S0(n8952), .S1(n8416), .Y(n8479) );
  MX4X1 U11848 ( .A(\buff[40][0] ), .B(\buff[44][0] ), .C(\buff[42][0] ), .D(
        \buff[46][0] ), .S0(n8952), .S1(n8416), .Y(n8478) );
  MXI2X1 U11849 ( .A(n8499), .B(n8498), .S0(n8923), .Y(n8747) );
  MX4X1 U11850 ( .A(\buff[8][1] ), .B(\buff[12][1] ), .C(\buff[10][1] ), .D(
        \buff[14][1] ), .S0(n8952), .S1(n8416), .Y(n8499) );
  MX4X1 U11851 ( .A(\buff[40][1] ), .B(\buff[44][1] ), .C(\buff[42][1] ), .D(
        \buff[46][1] ), .S0(n8952), .S1(n9152), .Y(n8498) );
  MXI2X1 U11852 ( .A(n8519), .B(n8518), .S0(n8923), .Y(n8754) );
  OAI21XL U11853 ( .A0(n621), .A1(n622), .B0(n623), .Y(n619) );
  OAI222XL U11854 ( .A0(n9420), .A1(n9602), .B0(n9356), .B1(n9421), .C0(n9599), 
        .C1(n9532), .Y(n622) );
  OAI21XL U11855 ( .A0(n630), .A1(n631), .B0(n623), .Y(n628) );
  OAI222XL U11856 ( .A0(n9420), .A1(n9592), .B0(n9355), .B1(n9421), .C0(n9588), 
        .C1(n9532), .Y(n631) );
  OAI21XL U11857 ( .A0(n635), .A1(n636), .B0(n623), .Y(n633) );
  OAI222XL U11858 ( .A0(n9420), .A1(n9583), .B0(n9354), .B1(n9421), .C0(n9581), 
        .C1(n9532), .Y(n636) );
  OAI21XL U11859 ( .A0(n640), .A1(n641), .B0(n623), .Y(n638) );
  OAI222XL U11860 ( .A0(n9420), .A1(n9574), .B0(n9353), .B1(n9421), .C0(n9572), 
        .C1(n9532), .Y(n641) );
  OAI21XL U11861 ( .A0(n645), .A1(n646), .B0(n623), .Y(n643) );
  OAI222XL U11862 ( .A0(n9420), .A1(n9564), .B0(n9352), .B1(n9421), .C0(n9563), 
        .C1(n9532), .Y(n646) );
  OAI21XL U11863 ( .A0(n650), .A1(n651), .B0(n623), .Y(n648) );
  OAI222XL U11864 ( .A0(n9420), .A1(n9557), .B0(n9351), .B1(n9421), .C0(n9554), 
        .C1(n9532), .Y(n651) );
  OAI21XL U11865 ( .A0(n655), .A1(n656), .B0(n623), .Y(n653) );
  OAI222XL U11866 ( .A0(n9420), .A1(n9546), .B0(n9350), .B1(n9421), .C0(n9545), 
        .C1(n9532), .Y(n656) );
  OAI21XL U11867 ( .A0(n660), .A1(n661), .B0(n623), .Y(n658) );
  OAI222XL U11868 ( .A0(n9420), .A1(n9537), .B0(n9346), .B1(n9421), .C0(n9536), 
        .C1(n9532), .Y(n661) );
  OAI21XL U11869 ( .A0(n1266), .A1(n1267), .B0(n1268), .Y(n1264) );
  OAI222XL U11870 ( .A0(n9602), .A1(n9400), .B0(n9356), .B1(n9531), .C0(n9598), 
        .C1(n9526), .Y(n1267) );
  OAI21XL U11871 ( .A0(n1274), .A1(n1275), .B0(n1268), .Y(n1272) );
  OAI222XL U11872 ( .A0(n320), .A1(n9400), .B0(n9355), .B1(n9531), .C0(n9589), 
        .C1(n9526), .Y(n1275) );
  OAI21XL U11873 ( .A0(n1278), .A1(n1279), .B0(n1268), .Y(n1276) );
  OAI222XL U11874 ( .A0(n9582), .A1(n9400), .B0(n9354), .B1(n9531), .C0(n9580), 
        .C1(n9526), .Y(n1279) );
  OAI21XL U11875 ( .A0(n1282), .A1(n1283), .B0(n1268), .Y(n1280) );
  OAI222XL U11876 ( .A0(n9573), .A1(n9400), .B0(n9353), .B1(n9531), .C0(n9571), 
        .C1(n9526), .Y(n1283) );
  OAI21XL U11877 ( .A0(n1286), .A1(n1287), .B0(n1268), .Y(n1284) );
  OAI222XL U11878 ( .A0(n9564), .A1(n9400), .B0(n9352), .B1(n9531), .C0(n345), 
        .C1(n9526), .Y(n1287) );
  OAI21XL U11879 ( .A0(n1290), .A1(n1291), .B0(n1268), .Y(n1288) );
  OAI222XL U11880 ( .A0(n9557), .A1(n9400), .B0(n9351), .B1(n9531), .C0(n9553), 
        .C1(n9526), .Y(n1291) );
  OAI21XL U11881 ( .A0(n1294), .A1(n1295), .B0(n1268), .Y(n1292) );
  OAI222XL U11882 ( .A0(n9548), .A1(n9400), .B0(n9350), .B1(n9531), .C0(n9544), 
        .C1(n9526), .Y(n1295) );
  OAI21XL U11883 ( .A0(n1298), .A1(n1299), .B0(n1268), .Y(n1296) );
  OAI222XL U11884 ( .A0(n9539), .A1(n9400), .B0(n9346), .B1(n9531), .C0(n9535), 
        .C1(n9526), .Y(n1299) );
  OAI21XL U11885 ( .A0(n1583), .A1(n1584), .B0(n1585), .Y(n1581) );
  OAI222XL U11886 ( .A0(n9601), .A1(n9390), .B0(n9356), .B1(n9527), .C0(n9598), 
        .C1(n9524), .Y(n1584) );
  OAI21XL U11887 ( .A0(n1591), .A1(n1592), .B0(n1585), .Y(n1589) );
  OAI222XL U11888 ( .A0(n9593), .A1(n9390), .B0(n9355), .B1(n9527), .C0(n9589), 
        .C1(n9524), .Y(n1592) );
  OAI21XL U11889 ( .A0(n1595), .A1(n1596), .B0(n1585), .Y(n1593) );
  OAI222XL U11890 ( .A0(n9582), .A1(n9390), .B0(n9354), .B1(n9527), .C0(n9580), 
        .C1(n9524), .Y(n1596) );
  OAI21XL U11891 ( .A0(n1599), .A1(n1600), .B0(n1585), .Y(n1597) );
  OAI222XL U11892 ( .A0(n9575), .A1(n9390), .B0(n9353), .B1(n9527), .C0(n9571), 
        .C1(n9524), .Y(n1600) );
  OAI21XL U11893 ( .A0(n1603), .A1(n1604), .B0(n1585), .Y(n1601) );
  OAI222XL U11894 ( .A0(n9566), .A1(n9390), .B0(n9352), .B1(n9527), .C0(n9561), 
        .C1(n9524), .Y(n1604) );
  OAI21XL U11895 ( .A0(n1607), .A1(n1608), .B0(n1585), .Y(n1605) );
  OAI222XL U11896 ( .A0(n9556), .A1(n9390), .B0(n9351), .B1(n9527), .C0(n9553), 
        .C1(n9524), .Y(n1608) );
  OAI21XL U11897 ( .A0(n1611), .A1(n1612), .B0(n1585), .Y(n1609) );
  OAI222XL U11898 ( .A0(n9548), .A1(n9390), .B0(n9350), .B1(n9527), .C0(n9544), 
        .C1(n9524), .Y(n1612) );
  OAI21XL U11899 ( .A0(n1615), .A1(n1616), .B0(n1585), .Y(n1613) );
  OAI222XL U11900 ( .A0(n9537), .A1(n9390), .B0(n9346), .B1(n9527), .C0(n9535), 
        .C1(n9524), .Y(n1616) );
  OAI21XL U11901 ( .A0(n1898), .A1(n1899), .B0(n1900), .Y(n1896) );
  OAI222XL U11902 ( .A0(n9600), .A1(n9523), .B0(n9356), .B1(n9525), .C0(n9597), 
        .C1(n9520), .Y(n1899) );
  OAI21XL U11903 ( .A0(n1906), .A1(n1907), .B0(n1900), .Y(n1904) );
  OAI222XL U11904 ( .A0(n9593), .A1(n9522), .B0(n9355), .B1(n9525), .C0(n9588), 
        .C1(n9520), .Y(n1907) );
  OAI21XL U11905 ( .A0(n1910), .A1(n1911), .B0(n1900), .Y(n1908) );
  OAI222XL U11906 ( .A0(n9584), .A1(n9522), .B0(n9354), .B1(n9525), .C0(n9579), 
        .C1(n9520), .Y(n1911) );
  OAI21XL U11907 ( .A0(n1914), .A1(n1915), .B0(n1900), .Y(n1912) );
  OAI222XL U11908 ( .A0(n9575), .A1(n9522), .B0(n9353), .B1(n9525), .C0(n9570), 
        .C1(n9520), .Y(n1915) );
  OAI21XL U11909 ( .A0(n1918), .A1(n1919), .B0(n1900), .Y(n1916) );
  OAI222XL U11910 ( .A0(n9565), .A1(n9522), .B0(n9352), .B1(n9525), .C0(n9562), 
        .C1(n9520), .Y(n1919) );
  OAI21XL U11911 ( .A0(n1922), .A1(n1923), .B0(n1900), .Y(n1920) );
  OAI222XL U11912 ( .A0(n9555), .A1(n9522), .B0(n9351), .B1(n9525), .C0(n9552), 
        .C1(n9520), .Y(n1923) );
  OAI21XL U11913 ( .A0(n1926), .A1(n1927), .B0(n1900), .Y(n1924) );
  OAI222XL U11914 ( .A0(n9547), .A1(n9522), .B0(n9350), .B1(n9525), .C0(n9543), 
        .C1(n9520), .Y(n1927) );
  OAI21XL U11915 ( .A0(n1930), .A1(n1931), .B0(n1900), .Y(n1928) );
  OAI222XL U11916 ( .A0(n9538), .A1(n9522), .B0(n9346), .B1(n9525), .C0(n9534), 
        .C1(n9520), .Y(n1931) );
  OAI21XL U11917 ( .A0(n2217), .A1(n2218), .B0(n2219), .Y(n2215) );
  OAI222XL U11918 ( .A0(n9600), .A1(n9371), .B0(n9356), .B1(n9521), .C0(n9597), 
        .C1(n7236), .Y(n2218) );
  OAI21XL U11919 ( .A0(n2225), .A1(n2226), .B0(n2219), .Y(n2223) );
  OAI222XL U11920 ( .A0(n9593), .A1(n9371), .B0(n9355), .B1(n9521), .C0(n9588), 
        .C1(n7236), .Y(n2226) );
  OAI21XL U11921 ( .A0(n2229), .A1(n2230), .B0(n2219), .Y(n2227) );
  OAI222XL U11922 ( .A0(n9584), .A1(n9371), .B0(n9354), .B1(n9521), .C0(n9579), 
        .C1(n7236), .Y(n2230) );
  OAI21XL U11923 ( .A0(n2233), .A1(n2234), .B0(n2219), .Y(n2231) );
  OAI222XL U11924 ( .A0(n9575), .A1(n9371), .B0(n9353), .B1(n9521), .C0(n9570), 
        .C1(n7236), .Y(n2234) );
  OAI21XL U11925 ( .A0(n2237), .A1(n2238), .B0(n2219), .Y(n2235) );
  OAI222XL U11926 ( .A0(n9565), .A1(n9371), .B0(n9352), .B1(n9521), .C0(n9562), 
        .C1(n7236), .Y(n2238) );
  OAI21XL U11927 ( .A0(n2241), .A1(n2242), .B0(n2219), .Y(n2239) );
  OAI222XL U11928 ( .A0(n9555), .A1(n9371), .B0(n9351), .B1(n9521), .C0(n9552), 
        .C1(n7236), .Y(n2242) );
  OAI21XL U11929 ( .A0(n2245), .A1(n2246), .B0(n2219), .Y(n2243) );
  OAI222XL U11930 ( .A0(n9547), .A1(n9371), .B0(n9350), .B1(n9521), .C0(n9543), 
        .C1(n7236), .Y(n2246) );
  OAI21XL U11931 ( .A0(n2249), .A1(n2250), .B0(n2219), .Y(n2247) );
  OAI222XL U11932 ( .A0(n9538), .A1(n9371), .B0(n9346), .B1(n9521), .C0(n9534), 
        .C1(n7236), .Y(n2250) );
  OAI21XL U11933 ( .A0(n962), .A1(n963), .B0(n948), .Y(n960) );
  OAI222XL U11934 ( .A0(n9573), .A1(n9410), .B0(n9353), .B1(n9533), .C0(n9572), 
        .C1(n9530), .Y(n963) );
  OAI21XL U11935 ( .A0(n966), .A1(n967), .B0(n948), .Y(n964) );
  OAI222XL U11936 ( .A0(n9564), .A1(n9410), .B0(n9352), .B1(n9533), .C0(n9563), 
        .C1(n9530), .Y(n967) );
  OAI21XL U11937 ( .A0(n970), .A1(n971), .B0(n948), .Y(n968) );
  OAI222XL U11938 ( .A0(n9557), .A1(n9410), .B0(n9351), .B1(n9533), .C0(n9554), 
        .C1(n9530), .Y(n971) );
  OAI21XL U11939 ( .A0(n974), .A1(n975), .B0(n948), .Y(n972) );
  OAI222XL U11940 ( .A0(n9548), .A1(n9410), .B0(n9350), .B1(n9533), .C0(n9545), 
        .C1(n9530), .Y(n975) );
  OAI21XL U11941 ( .A0(n978), .A1(n979), .B0(n948), .Y(n976) );
  OAI222XL U11942 ( .A0(n9539), .A1(n9410), .B0(n9346), .B1(n9533), .C0(n9536), 
        .C1(n9530), .Y(n979) );
  OAI21XL U11943 ( .A0(n1440), .A1(n1441), .B0(n1426), .Y(n1438) );
  OAI222XL U11944 ( .A0(n9573), .A1(n9396), .B0(n9353), .B1(n9529), .C0(n9571), 
        .C1(n9387), .Y(n1441) );
  OAI21XL U11945 ( .A0(n1444), .A1(n1445), .B0(n1426), .Y(n1442) );
  OAI222XL U11946 ( .A0(n9566), .A1(n9396), .B0(n9352), .B1(n9529), .C0(n345), 
        .C1(n9387), .Y(n1445) );
  OAI21XL U11947 ( .A0(n1448), .A1(n1449), .B0(n1426), .Y(n1446) );
  OAI222XL U11948 ( .A0(n9556), .A1(n9396), .B0(n9351), .B1(n9529), .C0(n9553), 
        .C1(n9387), .Y(n1449) );
  OAI21XL U11949 ( .A0(n1452), .A1(n1453), .B0(n1426), .Y(n1450) );
  OAI222XL U11950 ( .A0(n360), .A1(n9396), .B0(n9350), .B1(n9529), .C0(n9544), 
        .C1(n9387), .Y(n1453) );
  OAI21XL U11951 ( .A0(n1456), .A1(n1457), .B0(n1426), .Y(n1454) );
  OAI222XL U11952 ( .A0(n9539), .A1(n9396), .B0(n9346), .B1(n9529), .C0(n9535), 
        .C1(n9387), .Y(n1457) );
  OAI21XL U11953 ( .A0(n1953), .A1(n1954), .B0(n1939), .Y(n1951) );
  OAI222XL U11954 ( .A0(n9575), .A1(n9381), .B0(n9353), .B1(n9523), .C0(n9570), 
        .C1(n9371), .Y(n1954) );
  OAI21XL U11955 ( .A0(n1957), .A1(n1958), .B0(n1939), .Y(n1955) );
  OAI222XL U11956 ( .A0(n9565), .A1(n9381), .B0(n9352), .B1(n9523), .C0(n9562), 
        .C1(n9371), .Y(n1958) );
  OAI21XL U11957 ( .A0(n1961), .A1(n1962), .B0(n1939), .Y(n1959) );
  OAI222XL U11958 ( .A0(n9555), .A1(n9381), .B0(n9351), .B1(n9523), .C0(n9552), 
        .C1(n9371), .Y(n1962) );
  OAI21XL U11959 ( .A0(n1965), .A1(n1966), .B0(n1939), .Y(n1963) );
  OAI222XL U11960 ( .A0(n9547), .A1(n9381), .B0(n9350), .B1(n9523), .C0(n9543), 
        .C1(n9371), .Y(n1966) );
  OAI21XL U11961 ( .A0(n1969), .A1(n1970), .B0(n1939), .Y(n1967) );
  OAI222XL U11962 ( .A0(n9538), .A1(n9381), .B0(n9346), .B1(n9523), .C0(n9534), 
        .C1(n9371), .Y(n1970) );
  OAI21XL U11963 ( .A0(n2438), .A1(n2439), .B0(n2420), .Y(n2436) );
  OAI222XL U11964 ( .A0(n9561), .A1(n9361), .B0(n9352), .B1(n9519), .C0(n9564), 
        .C1(n9358), .Y(n2439) );
  OAI21XL U11965 ( .A0(n2442), .A1(n2443), .B0(n2420), .Y(n2440) );
  OAI222XL U11966 ( .A0(n9554), .A1(n9361), .B0(n9351), .B1(n9519), .C0(n9555), 
        .C1(n9358), .Y(n2443) );
  OAI21XL U11967 ( .A0(n2446), .A1(n2447), .B0(n2420), .Y(n2444) );
  OAI222XL U11968 ( .A0(n9545), .A1(n9361), .B0(n9350), .B1(n9519), .C0(n9546), 
        .C1(n9358), .Y(n2447) );
  OAI21XL U11969 ( .A0(n2450), .A1(n2451), .B0(n2420), .Y(n2448) );
  OAI222XL U11970 ( .A0(n9536), .A1(n9361), .B0(n9346), .B1(n9519), .C0(n9537), 
        .C1(n9358), .Y(n2451) );
  CLKMX2X2 U11971 ( .A(n8450), .B(n8451), .S0(n8922), .Y(n8492) );
  MX3XL U11972 ( .A(n8871), .B(n8863), .C(n8489), .S0(n8941), .S1(n8957), .Y(
        n8450) );
  MX3XL U11973 ( .A(n8823), .B(n8815), .C(n8488), .S0(n8942), .S1(n8957), .Y(
        n8451) );
  CLKMX2X2 U11974 ( .A(n8452), .B(n8453), .S0(n8923), .Y(n8512) );
  MX3XL U11975 ( .A(n8872), .B(n8864), .C(n8509), .S0(n8942), .S1(n8958), .Y(
        n8452) );
  MX3XL U11976 ( .A(n8824), .B(n8816), .C(n8508), .S0(n8942), .S1(n8958), .Y(
        n8453) );
  MXI2X1 U11977 ( .A(\buff[41][2] ), .B(\buff[45][2] ), .S0(n8431), .Y(n8528)
         );
  MXI2X1 U11978 ( .A(\buff[9][2] ), .B(\buff[13][2] ), .S0(n9141), .Y(n8529)
         );
  MXI3X1 U11979 ( .A(\buff[23][2] ), .B(\buff[27][2] ), .C(n8889), .S0(n8941), 
        .S1(n8958), .Y(n8531) );
  CLKINVX1 U11980 ( .A(n8670), .Y(n8889) );
  MXI2X1 U11981 ( .A(\buff[27][0] ), .B(\buff[31][0] ), .S0(n8944), .Y(n8645)
         );
  MXI2X1 U11982 ( .A(n8456), .B(n8738), .S0(n8922), .Y(n8741) );
  MX4X1 U11983 ( .A(\buff[56][0] ), .B(\buff[60][0] ), .C(\buff[58][0] ), .D(
        \buff[62][0] ), .S0(n8949), .S1(n8960), .Y(n8738) );
  MXI2X1 U11984 ( .A(n8457), .B(n8745), .S0(n8921), .Y(n8748) );
  MX4X1 U11985 ( .A(\buff[56][1] ), .B(\buff[60][1] ), .C(\buff[58][1] ), .D(
        \buff[62][1] ), .S0(n8949), .S1(n8960), .Y(n8745) );
  NOR2X1 U11986 ( .A(n982), .B(reset), .Y(n2412) );
  AND2X2 U11987 ( .A(n2412), .B(n2585), .Y(n2132) );
  OAI21XL U11988 ( .A0(n9440), .A1(n9439), .B0(n9668), .Y(n115) );
  OAI21XL U11989 ( .A0(n9438), .A1(n9437), .B0(n9668), .Y(n118) );
  MXI2X1 U11990 ( .A(n8492), .B(n8744), .S0(n9513), .Y(n8743) );
  MXI2X1 U11991 ( .A(n8895), .B(n8742), .S0(n8922), .Y(n8744) );
  CLKINVX1 U11992 ( .A(n8491), .Y(n8895) );
  MXI2X1 U11993 ( .A(n8512), .B(n8751), .S0(n9513), .Y(n8750) );
  MXI2X1 U11994 ( .A(n8896), .B(n8749), .S0(n8921), .Y(n8751) );
  CLKINVX1 U11995 ( .A(n8511), .Y(n8896) );
  MXI2X1 U11996 ( .A(n8532), .B(n8758), .S0(n8927), .Y(n8757) );
  MXI2X1 U11997 ( .A(n8897), .B(n8756), .S0(n9515), .Y(n8758) );
  MX4X1 U11998 ( .A(\buff[55][2] ), .B(\buff[59][2] ), .C(\buff[57][2] ), .D(
        \buff[61][2] ), .S0(n8948), .S1(n8960), .Y(n8756) );
  CLKINVX1 U11999 ( .A(n8531), .Y(n8897) );
  OAI2BB2XL U12000 ( .B0(n9432), .B1(n232), .A0N(\buff[55][0] ), .A1N(n9432), 
        .Y(n2658) );
  OAI222XL U12001 ( .A0(n9812), .A1(n238), .B0(n9725), .B1(n9431), .C0(n241), 
        .C1(n9804), .Y(n234) );
  OAI2BB2XL U12002 ( .B0(n9432), .B1(n243), .A0N(\buff[55][1] ), .A1N(n9432), 
        .Y(n2659) );
  OAI222XL U12003 ( .A0(n9811), .A1(n238), .B0(n9724), .B1(n9431), .C0(n241), 
        .C1(n9803), .Y(n244) );
  OAI2BB2XL U12004 ( .B0(n9432), .B1(n250), .A0N(\buff[55][2] ), .A1N(n9432), 
        .Y(n2660) );
  AOI211X1 U12005 ( .A0(n233), .A1(n8434), .B0(n251), .C0(n9446), .Y(n250) );
  OAI222XL U12006 ( .A0(n9810), .A1(n238), .B0(n9723), .B1(n9431), .C0(n241), 
        .C1(n9802), .Y(n251) );
  CLKINVX1 U12007 ( .A(n8434), .Y(n9802) );
  OAI2BB2XL U12008 ( .B0(n9432), .B1(n257), .A0N(\buff[55][3] ), .A1N(n9432), 
        .Y(n2661) );
  AOI211X1 U12009 ( .A0(n233), .A1(n8435), .B0(n258), .C0(n9444), .Y(n257) );
  OAI222XL U12010 ( .A0(n9809), .A1(n238), .B0(n9722), .B1(n9431), .C0(n241), 
        .C1(n9801), .Y(n258) );
  CLKINVX1 U12011 ( .A(n8435), .Y(n9801) );
  OAI2BB2XL U12012 ( .B0(n9432), .B1(n264), .A0N(n7446), .A1N(n9432), .Y(n2662) );
  AOI211X1 U12013 ( .A0(n233), .A1(n8442), .B0(n265), .C0(n9442), .Y(n264) );
  OAI222XL U12014 ( .A0(n9494), .A1(n238), .B0(n9721), .B1(n9431), .C0(n241), 
        .C1(n9800), .Y(n265) );
  CLKINVX1 U12015 ( .A(n8442), .Y(n9800) );
  OAI2BB2XL U12016 ( .B0(n9432), .B1(n271), .A0N(n7448), .A1N(n9432), .Y(n2663) );
  AOI211X1 U12017 ( .A0(n233), .A1(n8443), .B0(n272), .C0(n9440), .Y(n271) );
  OAI222XL U12018 ( .A0(n9491), .A1(n238), .B0(n9720), .B1(n9431), .C0(n241), 
        .C1(n9799), .Y(n272) );
  CLKINVX1 U12019 ( .A(n8443), .Y(n9799) );
  OAI2BB2XL U12020 ( .B0(n9432), .B1(n278), .A0N(n7528), .A1N(n9432), .Y(n2664) );
  AOI211X1 U12021 ( .A0(n233), .A1(n8444), .B0(n279), .C0(n9438), .Y(n278) );
  OAI222XL U12022 ( .A0(n9489), .A1(n238), .B0(n9719), .B1(n9431), .C0(n241), 
        .C1(n9798), .Y(n279) );
  CLKINVX1 U12023 ( .A(n8444), .Y(n9798) );
  OAI2BB2XL U12024 ( .B0(n9432), .B1(n285), .A0N(n7530), .A1N(n9432), .Y(n2665) );
  AOI211X1 U12025 ( .A0(n233), .A1(n8445), .B0(n286), .C0(n9436), .Y(n285) );
  OAI222XL U12026 ( .A0(n241), .A1(n9797), .B0(n9486), .B1(n238), .C0(n9718), 
        .C1(n9431), .Y(n286) );
  CLKINVX1 U12027 ( .A(n8445), .Y(n9797) );
  OAI2BB2XL U12028 ( .B0(n9456), .B1(n149), .A0N(\buff[61][0] ), .A1N(n9456), 
        .Y(n2610) );
  AOI221XL U12029 ( .A0(n9795), .A1(n128), .B0(n9429), .B1(n9449), .C0(n9450), 
        .Y(n149) );
  OAI2BB2XL U12030 ( .B0(n9456), .B1(n152), .A0N(\buff[61][1] ), .A1N(n9456), 
        .Y(n2611) );
  AOI221XL U12031 ( .A0(n9795), .A1(n131), .B0(n9429), .B1(n9447), .C0(n9448), 
        .Y(n152) );
  OAI2BB2XL U12032 ( .B0(n9456), .B1(n153), .A0N(\buff[61][2] ), .A1N(n9456), 
        .Y(n2612) );
  AOI221XL U12033 ( .A0(n9795), .A1(n133), .B0(n9429), .B1(n9445), .C0(n9446), 
        .Y(n153) );
  OAI2BB2XL U12034 ( .B0(n9456), .B1(n154), .A0N(\buff[61][3] ), .A1N(n9456), 
        .Y(n2613) );
  AOI221XL U12035 ( .A0(n9795), .A1(n135), .B0(n9429), .B1(n9443), .C0(n9444), 
        .Y(n154) );
  OAI2BB2XL U12036 ( .B0(n9456), .B1(n155), .A0N(n7313), .A1N(n9456), .Y(n2614) );
  AOI221XL U12037 ( .A0(n9795), .A1(n137), .B0(n9429), .B1(n9441), .C0(n9442), 
        .Y(n155) );
  OAI2BB2XL U12038 ( .B0(n9455), .B1(n163), .A0N(\buff[60][0] ), .A1N(n9455), 
        .Y(n2618) );
  AOI221XL U12039 ( .A0(n9794), .A1(n128), .B0(n9428), .B1(n9449), .C0(n9450), 
        .Y(n163) );
  OAI2BB2XL U12040 ( .B0(n9455), .B1(n166), .A0N(\buff[60][1] ), .A1N(n9455), 
        .Y(n2619) );
  AOI221XL U12041 ( .A0(n9794), .A1(n131), .B0(n9428), .B1(n9447), .C0(n9448), 
        .Y(n166) );
  OAI2BB2XL U12042 ( .B0(n9455), .B1(n167), .A0N(\buff[60][2] ), .A1N(n9455), 
        .Y(n2620) );
  AOI221XL U12043 ( .A0(n9794), .A1(n133), .B0(n9428), .B1(n9445), .C0(n9446), 
        .Y(n167) );
  OAI2BB2XL U12044 ( .B0(n9455), .B1(n168), .A0N(\buff[60][3] ), .A1N(n9455), 
        .Y(n2621) );
  AOI221XL U12045 ( .A0(n9794), .A1(n135), .B0(n9428), .B1(n9443), .C0(n9444), 
        .Y(n168) );
  OAI2BB2XL U12046 ( .B0(n9455), .B1(n169), .A0N(n7337), .A1N(n9455), .Y(n2622) );
  AOI221XL U12047 ( .A0(n9794), .A1(n137), .B0(n9428), .B1(n9441), .C0(n9442), 
        .Y(n169) );
  OAI2BB2XL U12048 ( .B0(n9454), .B1(n176), .A0N(\buff[59][0] ), .A1N(n9454), 
        .Y(n2626) );
  AOI221XL U12049 ( .A0(n9793), .A1(n128), .B0(n9427), .B1(n9449), .C0(n9450), 
        .Y(n176) );
  OAI2BB2XL U12050 ( .B0(n9454), .B1(n179), .A0N(\buff[59][1] ), .A1N(n9454), 
        .Y(n2627) );
  AOI221XL U12051 ( .A0(n9793), .A1(n131), .B0(n9427), .B1(n9447), .C0(n9448), 
        .Y(n179) );
  OAI2BB2XL U12052 ( .B0(n9454), .B1(n180), .A0N(\buff[59][2] ), .A1N(n9454), 
        .Y(n2628) );
  AOI221XL U12053 ( .A0(n9793), .A1(n133), .B0(n9427), .B1(n9445), .C0(n9446), 
        .Y(n180) );
  OAI2BB2XL U12054 ( .B0(n9454), .B1(n181), .A0N(\buff[59][3] ), .A1N(n9454), 
        .Y(n2629) );
  AOI221XL U12055 ( .A0(n9793), .A1(n135), .B0(n9427), .B1(n9443), .C0(n9444), 
        .Y(n181) );
  OAI2BB2XL U12056 ( .B0(n9454), .B1(n182), .A0N(n7360), .A1N(n9454), .Y(n2630) );
  AOI221XL U12057 ( .A0(n9793), .A1(n137), .B0(n9427), .B1(n9441), .C0(n9442), 
        .Y(n182) );
  OAI2BB2XL U12058 ( .B0(n9453), .B1(n189), .A0N(\buff[58][0] ), .A1N(n9453), 
        .Y(n2634) );
  AOI221XL U12059 ( .A0(n9792), .A1(n128), .B0(n9426), .B1(n9449), .C0(n9450), 
        .Y(n189) );
  OAI2BB2XL U12060 ( .B0(n9453), .B1(n192), .A0N(\buff[58][1] ), .A1N(n9453), 
        .Y(n2635) );
  AOI221XL U12061 ( .A0(n9792), .A1(n131), .B0(n9426), .B1(n9447), .C0(n9448), 
        .Y(n192) );
  OAI2BB2XL U12062 ( .B0(n9453), .B1(n193), .A0N(\buff[58][2] ), .A1N(n9453), 
        .Y(n2636) );
  AOI221XL U12063 ( .A0(n9792), .A1(n133), .B0(n9426), .B1(n9445), .C0(n9446), 
        .Y(n193) );
  OAI2BB2XL U12064 ( .B0(n9453), .B1(n194), .A0N(\buff[58][3] ), .A1N(n9453), 
        .Y(n2637) );
  AOI221XL U12065 ( .A0(n9792), .A1(n135), .B0(n9426), .B1(n9443), .C0(n9444), 
        .Y(n194) );
  OAI2BB2XL U12066 ( .B0(n9453), .B1(n195), .A0N(n7383), .A1N(n9453), .Y(n2638) );
  AOI221XL U12067 ( .A0(n9792), .A1(n137), .B0(n9426), .B1(n9441), .C0(n9442), 
        .Y(n195) );
  OAI2BB2XL U12068 ( .B0(n9452), .B1(n202), .A0N(\buff[57][0] ), .A1N(n9452), 
        .Y(n2642) );
  AOI221XL U12069 ( .A0(n9791), .A1(n128), .B0(n9425), .B1(n9449), .C0(n9450), 
        .Y(n202) );
  OAI2BB2XL U12070 ( .B0(n9452), .B1(n205), .A0N(\buff[57][1] ), .A1N(n9452), 
        .Y(n2643) );
  AOI221XL U12071 ( .A0(n9791), .A1(n131), .B0(n9425), .B1(n9447), .C0(n9448), 
        .Y(n205) );
  OAI2BB2XL U12072 ( .B0(n9452), .B1(n206), .A0N(\buff[57][2] ), .A1N(n9452), 
        .Y(n2644) );
  AOI221XL U12073 ( .A0(n9791), .A1(n133), .B0(n9425), .B1(n9445), .C0(n9446), 
        .Y(n206) );
  OAI2BB2XL U12074 ( .B0(n9452), .B1(n207), .A0N(\buff[57][3] ), .A1N(n9452), 
        .Y(n2645) );
  AOI221XL U12075 ( .A0(n9791), .A1(n135), .B0(n9425), .B1(n9443), .C0(n9444), 
        .Y(n207) );
  OAI2BB2XL U12076 ( .B0(n9452), .B1(n208), .A0N(n7407), .A1N(n9452), .Y(n2646) );
  AOI221XL U12077 ( .A0(n9791), .A1(n137), .B0(n9425), .B1(n9441), .C0(n9442), 
        .Y(n208) );
  OAI2BB2XL U12078 ( .B0(n9451), .B1(n215), .A0N(\buff[56][0] ), .A1N(n9451), 
        .Y(n2650) );
  AOI221XL U12079 ( .A0(n9790), .A1(n128), .B0(n9424), .B1(n9449), .C0(n9450), 
        .Y(n215) );
  OAI2BB2XL U12080 ( .B0(n9451), .B1(n220), .A0N(\buff[56][1] ), .A1N(n9451), 
        .Y(n2651) );
  AOI221XL U12081 ( .A0(n9790), .A1(n131), .B0(n9424), .B1(n9447), .C0(n9448), 
        .Y(n220) );
  OAI2BB2XL U12082 ( .B0(n9451), .B1(n221), .A0N(\buff[56][2] ), .A1N(n9451), 
        .Y(n2652) );
  AOI221XL U12083 ( .A0(n9790), .A1(n133), .B0(n9424), .B1(n9445), .C0(n9446), 
        .Y(n221) );
  OAI2BB2XL U12084 ( .B0(n9451), .B1(n222), .A0N(\buff[56][3] ), .A1N(n9451), 
        .Y(n2653) );
  AOI221XL U12085 ( .A0(n9790), .A1(n135), .B0(n9424), .B1(n9443), .C0(n9444), 
        .Y(n222) );
  OAI2BB2XL U12086 ( .B0(n9451), .B1(n223), .A0N(n7431), .A1N(n9451), .Y(n2654) );
  AOI221XL U12087 ( .A0(n9790), .A1(n137), .B0(n9424), .B1(n9441), .C0(n9442), 
        .Y(n223) );
  OAI2BB2XL U12088 ( .B0(n9457), .B1(n127), .A0N(\buff[62][0] ), .A1N(n9457), 
        .Y(n2602) );
  AOI221XL U12089 ( .A0(n9796), .A1(n128), .B0(n9449), .B1(n9430), .C0(n9450), 
        .Y(n127) );
  OAI2BB2XL U12090 ( .B0(n9457), .B1(n130), .A0N(\buff[62][1] ), .A1N(n9457), 
        .Y(n2603) );
  AOI221XL U12091 ( .A0(n9796), .A1(n131), .B0(n9447), .B1(n9430), .C0(n9448), 
        .Y(n130) );
  OAI2BB2XL U12092 ( .B0(n9457), .B1(n132), .A0N(\buff[62][2] ), .A1N(n9457), 
        .Y(n2604) );
  AOI221XL U12093 ( .A0(n9796), .A1(n133), .B0(n9445), .B1(n9430), .C0(n9446), 
        .Y(n132) );
  OAI2BB2XL U12094 ( .B0(n9457), .B1(n134), .A0N(\buff[62][3] ), .A1N(n9457), 
        .Y(n2605) );
  AOI221XL U12095 ( .A0(n9796), .A1(n135), .B0(n9443), .B1(n9430), .C0(n9444), 
        .Y(n134) );
  OAI2BB2XL U12096 ( .B0(n9457), .B1(n136), .A0N(n7289), .A1N(n9457), .Y(n2606) );
  AOI221XL U12097 ( .A0(n9796), .A1(n137), .B0(n9441), .B1(n9430), .C0(n9442), 
        .Y(n136) );
  CLKMX2X2 U12098 ( .A(n8454), .B(n8455), .S0(n8923), .Y(n8532) );
  MX3XL U12099 ( .A(n8873), .B(n8865), .C(n8529), .S0(n8942), .S1(n8958), .Y(
        n8454) );
  MX3XL U12100 ( .A(n8825), .B(n8817), .C(n8528), .S0(n8941), .S1(n8958), .Y(
        n8455) );
  MX4X1 U12101 ( .A(\buff[4][0] ), .B(\buff[5][0] ), .C(\buff[6][0] ), .D(
        \buff[7][0] ), .S0(n9134), .S1(n9147), .Y(n8982) );
  MX4X1 U12102 ( .A(\buff[36][0] ), .B(\buff[37][0] ), .C(\buff[38][0] ), .D(
        \buff[39][0] ), .S0(n9135), .S1(n9146), .Y(n8972) );
  MX4X1 U12103 ( .A(\buff[4][1] ), .B(\buff[5][1] ), .C(\buff[6][1] ), .D(
        \buff[7][1] ), .S0(n9133), .S1(n9148), .Y(n9002) );
  MX4X1 U12104 ( .A(\buff[36][1] ), .B(\buff[37][1] ), .C(\buff[38][1] ), .D(
        \buff[39][1] ), .S0(n9134), .S1(n9147), .Y(n8992) );
  MX4X1 U12105 ( .A(\buff[52][0] ), .B(\buff[53][0] ), .C(\buff[54][0] ), .D(
        \buff[55][0] ), .S0(n9135), .S1(n9146), .Y(n8967) );
  MX4X1 U12106 ( .A(n8978), .B(n8976), .C(n8977), .D(n8975), .S0(n9139), .S1(
        n9140), .Y(n8979) );
  MX4X1 U12107 ( .A(\buff[24][0] ), .B(\buff[25][0] ), .C(\buff[26][0] ), .D(
        \buff[27][0] ), .S0(n9135), .S1(n9146), .Y(n8976) );
  MX4X1 U12108 ( .A(\buff[28][0] ), .B(\buff[29][0] ), .C(\buff[30][0] ), .D(
        \buff[31][0] ), .S0(n9135), .S1(n9146), .Y(n8975) );
  MX4X1 U12109 ( .A(\buff[20][0] ), .B(\buff[21][0] ), .C(\buff[22][0] ), .D(
        \buff[23][0] ), .S0(n9135), .S1(n9146), .Y(n8977) );
  MX4X1 U12110 ( .A(\buff[20][1] ), .B(\buff[21][1] ), .C(\buff[22][1] ), .D(
        \buff[23][1] ), .S0(n9133), .S1(n9148), .Y(n8997) );
  MX4X1 U12111 ( .A(\buff[52][1] ), .B(\buff[53][1] ), .C(\buff[54][1] ), .D(
        \buff[55][1] ), .S0(n9134), .S1(n9147), .Y(n8987) );
  MX4X1 U12112 ( .A(n8998), .B(n8996), .C(n8997), .D(n8995), .S0(n9139), .S1(
        n8431), .Y(n8999) );
  MX4X1 U12113 ( .A(\buff[16][1] ), .B(\buff[17][1] ), .C(\buff[18][1] ), .D(
        \buff[19][1] ), .S0(n9133), .S1(n9148), .Y(n8998) );
  MX4X1 U12114 ( .A(\buff[24][1] ), .B(\buff[25][1] ), .C(\buff[26][1] ), .D(
        \buff[27][1] ), .S0(n9134), .S1(n9148), .Y(n8996) );
  MX4X1 U12115 ( .A(\buff[28][1] ), .B(\buff[29][1] ), .C(\buff[30][1] ), .D(
        \buff[31][1] ), .S0(n9134), .S1(n9148), .Y(n8995) );
  MX4X1 U12116 ( .A(\buff[16][0] ), .B(\buff[17][0] ), .C(\buff[18][0] ), .D(
        \buff[19][0] ), .S0(n9135), .S1(n9147), .Y(n8978) );
  MX4X1 U12117 ( .A(\buff[0][0] ), .B(\buff[1][0] ), .C(\buff[2][0] ), .D(
        \buff[3][0] ), .S0(n9134), .S1(n9147), .Y(n8983) );
  MX4X1 U12118 ( .A(\buff[48][0] ), .B(\buff[49][0] ), .C(\buff[50][0] ), .D(
        \buff[51][0] ), .S0(n9135), .S1(n9146), .Y(n8968) );
  MX4X1 U12119 ( .A(\buff[32][0] ), .B(\buff[33][0] ), .C(\buff[34][0] ), .D(
        \buff[35][0] ), .S0(n9135), .S1(n9146), .Y(n8973) );
  MX4X1 U12120 ( .A(\buff[48][1] ), .B(\buff[49][1] ), .C(\buff[50][1] ), .D(
        \buff[51][1] ), .S0(n9134), .S1(n9147), .Y(n8988) );
  MX4X1 U12121 ( .A(\buff[12][0] ), .B(\buff[13][0] ), .C(\buff[14][0] ), .D(
        \buff[15][0] ), .S0(n9135), .S1(n9147), .Y(n8980) );
  MX4X1 U12122 ( .A(\buff[44][0] ), .B(\buff[45][0] ), .C(\buff[46][0] ), .D(
        \buff[47][0] ), .S0(n9135), .S1(n9146), .Y(n8970) );
  MX4X1 U12123 ( .A(\buff[12][1] ), .B(\buff[13][1] ), .C(\buff[14][1] ), .D(
        \buff[15][1] ), .S0(n9133), .S1(n9148), .Y(n9000) );
  MX4X1 U12124 ( .A(\buff[44][1] ), .B(\buff[45][1] ), .C(\buff[46][1] ), .D(
        \buff[47][1] ), .S0(n9134), .S1(n9147), .Y(n8990) );
  MX4X1 U12125 ( .A(\buff[60][0] ), .B(\buff[61][0] ), .C(\buff[62][0] ), .D(
        \buff[63][0] ), .S0(n9135), .S1(n9146), .Y(n8965) );
  MX4X1 U12126 ( .A(\buff[60][1] ), .B(\buff[61][1] ), .C(\buff[62][1] ), .D(
        \buff[63][1] ), .S0(n9134), .S1(n9147), .Y(n8985) );
  MX4X1 U12127 ( .A(\buff[8][0] ), .B(\buff[9][0] ), .C(\buff[10][0] ), .D(
        \buff[11][0] ), .S0(n9134), .S1(n9147), .Y(n8981) );
  MX4X1 U12128 ( .A(\buff[40][0] ), .B(\buff[41][0] ), .C(\buff[42][0] ), .D(
        \buff[43][0] ), .S0(n9135), .S1(n9146), .Y(n8971) );
  MX4X1 U12129 ( .A(\buff[56][0] ), .B(\buff[57][0] ), .C(\buff[58][0] ), .D(
        \buff[59][0] ), .S0(n9135), .S1(n9146), .Y(n8966) );
  MX4X1 U12130 ( .A(\buff[56][1] ), .B(\buff[57][1] ), .C(\buff[58][1] ), .D(
        \buff[59][1] ), .S0(n9134), .S1(n9147), .Y(n8986) );
  MX4X1 U12131 ( .A(\buff[0][0] ), .B(\buff[4][0] ), .C(\buff[2][0] ), .D(
        \buff[6][0] ), .S0(n8952), .S1(n9152), .Y(n8477) );
  MX4X1 U12132 ( .A(\buff[16][0] ), .B(\buff[20][0] ), .C(\buff[18][0] ), .D(
        \buff[22][0] ), .S0(n8952), .S1(n9145), .Y(n8475) );
  CLKBUFX3 U12133 ( .A(n9814), .Y(n9508) );
  CLKINVX1 U12134 ( .A(n2576), .Y(n9814) );
  MXI3X1 U12135 ( .A(n8855), .B(n8847), .C(n8483), .S0(n8941), .S1(n8957), .Y(
        n8482) );
  CLKINVX1 U12136 ( .A(\buff[19][0] ), .Y(n8847) );
  CLKINVX1 U12137 ( .A(\buff[15][0] ), .Y(n8855) );
  MXI3X1 U12138 ( .A(n8856), .B(n8848), .C(n8503), .S0(n8942), .S1(n8958), .Y(
        n8502) );
  CLKINVX1 U12139 ( .A(\buff[15][1] ), .Y(n8856) );
  CLKINVX1 U12140 ( .A(\buff[19][1] ), .Y(n8848) );
  MXI3X1 U12141 ( .A(n8857), .B(n8849), .C(n8523), .S0(n8942), .S1(n8958), .Y(
        n8522) );
  CLKINVX1 U12142 ( .A(\buff[19][2] ), .Y(n8849) );
  CLKINVX1 U12143 ( .A(\buff[15][2] ), .Y(n8857) );
  MX4X1 U12144 ( .A(\buff[24][0] ), .B(\buff[28][0] ), .C(\buff[26][0] ), .D(
        \buff[30][0] ), .S0(n8940), .S1(n8960), .Y(n8456) );
  MX4X1 U12145 ( .A(\buff[24][1] ), .B(\buff[28][1] ), .C(\buff[26][1] ), .D(
        \buff[30][1] ), .S0(n8941), .S1(n8959), .Y(n8457) );
  MXI4X1 U12146 ( .A(n8489), .B(n8641), .C(n8488), .D(n8642), .S0(n8961), .S1(
        n8921), .Y(n8640) );
  MXI2X1 U12147 ( .A(\buff[43][0] ), .B(\buff[47][0] ), .S0(n8945), .Y(n8642)
         );
  MXI2X1 U12148 ( .A(\buff[11][0] ), .B(\buff[15][0] ), .S0(n8944), .Y(n8641)
         );
  MXI4X1 U12149 ( .A(n8509), .B(n8654), .C(n8508), .D(n8655), .S0(n8961), .S1(
        n8921), .Y(n8653) );
  MXI2X1 U12150 ( .A(\buff[43][1] ), .B(\buff[47][1] ), .S0(n8944), .Y(n8655)
         );
  MXI2X1 U12151 ( .A(\buff[11][1] ), .B(\buff[15][1] ), .S0(n8943), .Y(n8654)
         );
  MXI2X1 U12152 ( .A(\buff[51][0] ), .B(\buff[55][0] ), .S0(n8945), .Y(n8636)
         );
  MXI2X1 U12153 ( .A(\buff[19][0] ), .B(\buff[23][0] ), .S0(n8945), .Y(n8635)
         );
  MXI2X1 U12154 ( .A(\buff[51][1] ), .B(\buff[55][1] ), .S0(n8944), .Y(n8649)
         );
  MXI2X1 U12155 ( .A(\buff[19][1] ), .B(\buff[23][1] ), .S0(n8944), .Y(n8648)
         );
  MXI2X1 U12156 ( .A(\buff[35][0] ), .B(\buff[39][0] ), .S0(n8945), .Y(n8639)
         );
  MXI2X1 U12157 ( .A(\buff[3][0] ), .B(\buff[7][0] ), .S0(n8945), .Y(n8638) );
  MXI2X1 U12158 ( .A(\buff[35][1] ), .B(\buff[39][1] ), .S0(n8944), .Y(n8652)
         );
  MXI2X1 U12159 ( .A(\buff[3][1] ), .B(\buff[7][1] ), .S0(n8944), .Y(n8651) );
  OAI21XL U12160 ( .A0(n9450), .A1(n9449), .B0(n9668), .Y(n99) );
  OAI21XL U12161 ( .A0(n9448), .A1(n9447), .B0(n9668), .Y(n103) );
  OAI21XL U12162 ( .A0(n9446), .A1(n9445), .B0(n9668), .Y(n106) );
  OAI21XL U12163 ( .A0(n9444), .A1(n9443), .B0(n9668), .Y(n109) );
  OAI21XL U12164 ( .A0(n9442), .A1(n9441), .B0(n9668), .Y(n112) );
  OAI21XL U12165 ( .A0(n9436), .A1(n9435), .B0(n9668), .Y(n121) );
  MX4X1 U12166 ( .A(\buff[48][0] ), .B(\buff[52][0] ), .C(\buff[50][0] ), .D(
        \buff[54][0] ), .S0(n8952), .S1(n8956), .Y(n8474) );
  MX4X1 U12167 ( .A(\buff[32][0] ), .B(\buff[36][0] ), .C(\buff[34][0] ), .D(
        \buff[38][0] ), .S0(n8952), .S1(n9152), .Y(n8476) );
  MX4X1 U12168 ( .A(\buff[48][1] ), .B(\buff[52][1] ), .C(\buff[50][1] ), .D(
        \buff[54][1] ), .S0(n8952), .S1(n9152), .Y(n8494) );
  MX4X1 U12169 ( .A(\buff[32][1] ), .B(\buff[36][1] ), .C(\buff[34][1] ), .D(
        \buff[38][1] ), .S0(n8952), .S1(n9145), .Y(n8496) );
  MX4X1 U12170 ( .A(\buff[48][2] ), .B(\buff[52][2] ), .C(\buff[50][2] ), .D(
        \buff[54][2] ), .S0(n8952), .S1(n9144), .Y(n8514) );
  MX4X1 U12171 ( .A(\buff[32][2] ), .B(\buff[36][2] ), .C(\buff[34][2] ), .D(
        \buff[38][2] ), .S0(n8951), .S1(n9144), .Y(n8516) );
  MX4X1 U12172 ( .A(\buff[48][3] ), .B(\buff[52][3] ), .C(\buff[50][3] ), .D(
        \buff[54][3] ), .S0(n8951), .S1(n9142), .Y(n8534) );
  MX4X1 U12173 ( .A(\buff[32][3] ), .B(\buff[36][3] ), .C(\buff[34][3] ), .D(
        \buff[38][3] ), .S0(n8951), .S1(n9142), .Y(n8536) );
  MXI2X1 U12174 ( .A(\buff[25][3] ), .B(\buff[29][3] ), .S0(n8946), .Y(n8683)
         );
  MXI2X1 U12175 ( .A(\buff[25][4] ), .B(\buff[29][4] ), .S0(n8946), .Y(n8696)
         );
  MXI2X1 U12176 ( .A(\buff[25][5] ), .B(\buff[29][5] ), .S0(n8937), .Y(n8709)
         );
  MXI2X1 U12177 ( .A(\buff[25][6] ), .B(\buff[29][6] ), .S0(n8938), .Y(n8722)
         );
  MXI2X1 U12178 ( .A(\buff[25][7] ), .B(\buff[29][7] ), .S0(n8945), .Y(n8735)
         );
  MXI2X1 U12179 ( .A(n8539), .B(n8538), .S0(n8923), .Y(n8761) );
  MXI2X1 U12180 ( .A(n8559), .B(n8558), .S0(n8923), .Y(n8768) );
  MXI2X1 U12181 ( .A(n8579), .B(n8578), .S0(n8923), .Y(n8775) );
  MXI2X1 U12182 ( .A(n8599), .B(n8598), .S0(n9136), .Y(n8782) );
  MXI2X1 U12183 ( .A(n8619), .B(n8618), .S0(n8923), .Y(n8789) );
  MX4X1 U12184 ( .A(\buff[40][7] ), .B(\buff[44][7] ), .C(\buff[42][7] ), .D(
        \buff[46][7] ), .S0(n8949), .S1(n8960), .Y(n8618) );
  OAI21XL U12185 ( .A0(n946), .A1(n947), .B0(n948), .Y(n944) );
  OAI222XL U12186 ( .A0(n9602), .A1(n9410), .B0(n9356), .B1(n9533), .C0(n9599), 
        .C1(n9530), .Y(n947) );
  OAI21XL U12187 ( .A0(n954), .A1(n955), .B0(n948), .Y(n952) );
  OAI222XL U12188 ( .A0(n9593), .A1(n9410), .B0(n9355), .B1(n9533), .C0(n321), 
        .C1(n9530), .Y(n955) );
  OAI21XL U12189 ( .A0(n958), .A1(n959), .B0(n948), .Y(n956) );
  OAI222XL U12190 ( .A0(n9582), .A1(n9410), .B0(n9354), .B1(n9533), .C0(n9581), 
        .C1(n9530), .Y(n959) );
  OAI21XL U12191 ( .A0(n1424), .A1(n1425), .B0(n1426), .Y(n1422) );
  OAI222XL U12192 ( .A0(n9601), .A1(n9396), .B0(n9356), .B1(n9529), .C0(n9598), 
        .C1(n9387), .Y(n1425) );
  OAI21XL U12193 ( .A0(n1432), .A1(n1433), .B0(n1426), .Y(n1430) );
  OAI222XL U12194 ( .A0(n9591), .A1(n9396), .B0(n9355), .B1(n9529), .C0(n9589), 
        .C1(n9387), .Y(n1433) );
  OAI21XL U12195 ( .A0(n1436), .A1(n1437), .B0(n1426), .Y(n1434) );
  OAI222XL U12196 ( .A0(n9582), .A1(n9396), .B0(n9354), .B1(n9529), .C0(n9580), 
        .C1(n9387), .Y(n1437) );
  OAI21XL U12197 ( .A0(n1937), .A1(n1938), .B0(n1939), .Y(n1935) );
  OAI222XL U12198 ( .A0(n9600), .A1(n9381), .B0(n9356), .B1(n9523), .C0(n9597), 
        .C1(n9371), .Y(n1938) );
  OAI21XL U12199 ( .A0(n1945), .A1(n1946), .B0(n1939), .Y(n1943) );
  OAI222XL U12200 ( .A0(n9593), .A1(n9381), .B0(n9355), .B1(n9523), .C0(n9588), 
        .C1(n9371), .Y(n1946) );
  OAI21XL U12201 ( .A0(n1949), .A1(n1950), .B0(n1939), .Y(n1947) );
  OAI222XL U12202 ( .A0(n9584), .A1(n9381), .B0(n9354), .B1(n9523), .C0(n9579), 
        .C1(n9371), .Y(n1950) );
  OAI21XL U12203 ( .A0(n2418), .A1(n2419), .B0(n2420), .Y(n2416) );
  OAI222XL U12204 ( .A0(n313), .A1(n9361), .B0(n9356), .B1(n9519), .C0(n9602), 
        .C1(n9358), .Y(n2419) );
  OAI21XL U12205 ( .A0(n2426), .A1(n2427), .B0(n2420), .Y(n2424) );
  OAI222XL U12206 ( .A0(n9590), .A1(n9361), .B0(n9355), .B1(n9519), .C0(n9592), 
        .C1(n9358), .Y(n2427) );
  OAI21XL U12207 ( .A0(n2430), .A1(n2431), .B0(n2420), .Y(n2428) );
  OAI222XL U12208 ( .A0(n9580), .A1(n9361), .B0(n9354), .B1(n9519), .C0(n9583), 
        .C1(n9358), .Y(n2431) );
  OAI21XL U12209 ( .A0(n2434), .A1(n2435), .B0(n2420), .Y(n2432) );
  OAI222XL U12210 ( .A0(n9571), .A1(n9361), .B0(n9353), .B1(n9519), .C0(n9574), 
        .C1(n9358), .Y(n2435) );
  MXI2X1 U12211 ( .A(\buff[1][3] ), .B(\buff[5][3] ), .S0(n9141), .Y(n8547) );
  MXI2X1 U12212 ( .A(\buff[1][4] ), .B(\buff[5][4] ), .S0(n8946), .Y(n8567) );
  MXI2X1 U12213 ( .A(\buff[1][5] ), .B(\buff[5][5] ), .S0(n8937), .Y(n8587) );
  MXI2X1 U12214 ( .A(\buff[1][6] ), .B(\buff[5][6] ), .S0(n8939), .Y(n8607) );
  MXI2X1 U12215 ( .A(\buff[33][3] ), .B(\buff[37][3] ), .S0(n9140), .Y(n8545)
         );
  MXI2X1 U12216 ( .A(\buff[41][3] ), .B(\buff[45][3] ), .S0(n8431), .Y(n8548)
         );
  MXI2X1 U12217 ( .A(\buff[49][3] ), .B(\buff[53][3] ), .S0(n8431), .Y(n8541)
         );
  MXI2X1 U12218 ( .A(\buff[33][4] ), .B(\buff[37][4] ), .S0(n8946), .Y(n8565)
         );
  MXI2X1 U12219 ( .A(\buff[41][4] ), .B(\buff[45][4] ), .S0(n8946), .Y(n8568)
         );
  MXI2X1 U12220 ( .A(\buff[49][4] ), .B(\buff[53][4] ), .S0(n8946), .Y(n8561)
         );
  MXI2X1 U12221 ( .A(\buff[33][5] ), .B(\buff[37][5] ), .S0(n9140), .Y(n8585)
         );
  MXI2X1 U12222 ( .A(\buff[41][5] ), .B(\buff[45][5] ), .S0(n8944), .Y(n8588)
         );
  MXI2X1 U12223 ( .A(\buff[49][5] ), .B(\buff[53][5] ), .S0(n9140), .Y(n8581)
         );
  MXI2X1 U12224 ( .A(\buff[33][6] ), .B(\buff[37][6] ), .S0(n8942), .Y(n8605)
         );
  MXI2X1 U12225 ( .A(\buff[41][6] ), .B(\buff[45][6] ), .S0(n8950), .Y(n8608)
         );
  MXI2X1 U12226 ( .A(\buff[49][6] ), .B(\buff[53][6] ), .S0(n8950), .Y(n8601)
         );
  MXI2X1 U12227 ( .A(\buff[33][7] ), .B(\buff[37][7] ), .S0(n8945), .Y(n8625)
         );
  MXI2X1 U12228 ( .A(\buff[49][7] ), .B(\buff[53][7] ), .S0(n8945), .Y(n8621)
         );
  MXI2X1 U12229 ( .A(\buff[17][3] ), .B(\buff[21][3] ), .S0(n9141), .Y(n8543)
         );
  MXI2X1 U12230 ( .A(\buff[17][4] ), .B(\buff[21][4] ), .S0(n8946), .Y(n8563)
         );
  MXI2X1 U12231 ( .A(\buff[17][5] ), .B(\buff[21][5] ), .S0(n8937), .Y(n8583)
         );
  MXI2X1 U12232 ( .A(\buff[17][6] ), .B(\buff[21][6] ), .S0(n8943), .Y(n8603)
         );
  MXI2X1 U12233 ( .A(\buff[17][7] ), .B(\buff[21][7] ), .S0(n8945), .Y(n8623)
         );
  MXI2X1 U12234 ( .A(\buff[9][3] ), .B(\buff[13][3] ), .S0(n8946), .Y(n8549)
         );
  MXI2X1 U12235 ( .A(\buff[9][4] ), .B(\buff[13][4] ), .S0(n8946), .Y(n8569)
         );
  MXI2X1 U12236 ( .A(\buff[9][5] ), .B(\buff[13][5] ), .S0(n8942), .Y(n8589)
         );
  MXI2X1 U12237 ( .A(\buff[9][6] ), .B(\buff[13][6] ), .S0(n8941), .Y(n8609)
         );
  MXI3X1 U12238 ( .A(\buff[23][3] ), .B(\buff[27][3] ), .C(n8890), .S0(n8941), 
        .S1(n8958), .Y(n8551) );
  CLKINVX1 U12239 ( .A(n8683), .Y(n8890) );
  MXI3X1 U12240 ( .A(\buff[23][4] ), .B(\buff[27][4] ), .C(n8891), .S0(n8941), 
        .S1(n8957), .Y(n8571) );
  CLKINVX1 U12241 ( .A(n8696), .Y(n8891) );
  MXI3X1 U12242 ( .A(\buff[23][5] ), .B(\buff[27][5] ), .C(n8892), .S0(n8942), 
        .S1(n8957), .Y(n8591) );
  CLKINVX1 U12243 ( .A(n8709), .Y(n8892) );
  MXI3X1 U12244 ( .A(\buff[23][6] ), .B(\buff[27][6] ), .C(n8893), .S0(n8942), 
        .S1(n8957), .Y(n8611) );
  CLKINVX1 U12245 ( .A(n8722), .Y(n8893) );
  MXI3X1 U12246 ( .A(\buff[23][7] ), .B(\buff[27][7] ), .C(n8894), .S0(n8942), 
        .S1(n8957), .Y(n8631) );
  CLKINVX1 U12247 ( .A(n8735), .Y(n8894) );
  NOR3X1 U12248 ( .A(n9717), .B(reset), .C(n9664), .Y(n2593) );
  NAND2X1 U12249 ( .A(IROM_Q[0]), .B(n9744), .Y(n236) );
  NAND2X1 U12250 ( .A(IROM_Q[1]), .B(n9744), .Y(n246) );
  NAND2X1 U12251 ( .A(IROM_Q[2]), .B(n9744), .Y(n253) );
  NAND2X1 U12252 ( .A(IROM_Q[3]), .B(n9744), .Y(n260) );
  NAND2X1 U12253 ( .A(IROM_Q[4]), .B(n9744), .Y(n267) );
  NAND2X1 U12254 ( .A(IROM_Q[5]), .B(n9744), .Y(n274) );
  NAND2X1 U12255 ( .A(IROM_Q[6]), .B(n9744), .Y(n281) );
  NAND2X1 U12256 ( .A(IROM_Q[7]), .B(n9744), .Y(n288) );
  MXI2X1 U12257 ( .A(\buff[27][1] ), .B(\buff[31][1] ), .S0(n8943), .Y(n8658)
         );
  MXI2X1 U12258 ( .A(\buff[27][2] ), .B(\buff[31][2] ), .S0(n8953), .Y(n8671)
         );
  MXI2X1 U12259 ( .A(\buff[27][3] ), .B(\buff[31][3] ), .S0(n8943), .Y(n8684)
         );
  MXI2X1 U12260 ( .A(\buff[27][4] ), .B(\buff[31][4] ), .S0(n8944), .Y(n8697)
         );
  MXI2X1 U12261 ( .A(\buff[27][5] ), .B(\buff[31][5] ), .S0(n9140), .Y(n8710)
         );
  MXI2X1 U12262 ( .A(n8466), .B(n8752), .S0(n9515), .Y(n8755) );
  MXI2X1 U12263 ( .A(n8467), .B(n8759), .S0(n9136), .Y(n8762) );
  MX4X1 U12264 ( .A(\buff[56][3] ), .B(\buff[60][3] ), .C(\buff[58][3] ), .D(
        \buff[62][3] ), .S0(n8948), .S1(n8960), .Y(n8759) );
  MXI2X1 U12265 ( .A(n8468), .B(n8766), .S0(n9136), .Y(n8769) );
  MX4X1 U12266 ( .A(\buff[56][4] ), .B(\buff[60][4] ), .C(\buff[58][4] ), .D(
        \buff[62][4] ), .S0(n8948), .S1(n8960), .Y(n8766) );
  MXI2X1 U12267 ( .A(n8469), .B(n8773), .S0(n8921), .Y(n8776) );
  MXI2X1 U12268 ( .A(n8470), .B(n8780), .S0(n8921), .Y(n8783) );
  MX4X1 U12269 ( .A(\buff[56][6] ), .B(\buff[60][6] ), .C(\buff[58][6] ), .D(
        \buff[62][6] ), .S0(n8948), .S1(n8960), .Y(n8780) );
  OAI211X1 U12270 ( .A0(n92), .A1(n8372), .B0(n2559), .C0(n9663), .Y(n2560) );
  OAI221XL U12271 ( .A0(n9665), .A1(n9717), .B0(IRB_RW), .B1(n9746), .C0(n2562), .Y(n2559) );
  NOR2X1 U12272 ( .A(n96), .B(n985), .Y(n2562) );
  MXI2X1 U12273 ( .A(n8552), .B(n8765), .S0(n8927), .Y(n8764) );
  MXI2X1 U12274 ( .A(n8898), .B(n8763), .S0(n9136), .Y(n8765) );
  MX4X1 U12275 ( .A(\buff[55][3] ), .B(\buff[59][3] ), .C(\buff[57][3] ), .D(
        \buff[61][3] ), .S0(n8948), .S1(n8960), .Y(n8763) );
  CLKINVX1 U12276 ( .A(n8551), .Y(n8898) );
  MXI2X1 U12277 ( .A(n8572), .B(n8772), .S0(n9137), .Y(n8771) );
  MXI2X1 U12278 ( .A(n8899), .B(n8770), .S0(n8921), .Y(n8772) );
  MX4X1 U12279 ( .A(\buff[55][4] ), .B(\buff[59][4] ), .C(\buff[57][4] ), .D(
        \buff[61][4] ), .S0(n8948), .S1(n8960), .Y(n8770) );
  CLKINVX1 U12280 ( .A(n8571), .Y(n8899) );
  MXI2X1 U12281 ( .A(n8592), .B(n8779), .S0(n8927), .Y(n8778) );
  MXI2X1 U12282 ( .A(n8900), .B(n8777), .S0(n8921), .Y(n8779) );
  MX4X1 U12283 ( .A(\buff[55][5] ), .B(\buff[59][5] ), .C(\buff[57][5] ), .D(
        \buff[61][5] ), .S0(n8948), .S1(n8960), .Y(n8777) );
  CLKINVX1 U12284 ( .A(n8591), .Y(n8900) );
  MXI2X1 U12285 ( .A(n8612), .B(n8786), .S0(n8927), .Y(n8785) );
  MXI2X1 U12286 ( .A(n8901), .B(n8784), .S0(n8921), .Y(n8786) );
  MX4X1 U12287 ( .A(\buff[55][6] ), .B(\buff[59][6] ), .C(\buff[57][6] ), .D(
        \buff[61][6] ), .S0(n8948), .S1(n8960), .Y(n8784) );
  CLKINVX1 U12288 ( .A(n8611), .Y(n8901) );
  MXI2X1 U12289 ( .A(n8632), .B(n8793), .S0(n9513), .Y(n8792) );
  MXI2X1 U12290 ( .A(n8902), .B(n8791), .S0(n9136), .Y(n8793) );
  MX4X1 U12291 ( .A(\buff[55][7] ), .B(\buff[59][7] ), .C(\buff[57][7] ), .D(
        \buff[61][7] ), .S0(n8948), .S1(n8960), .Y(n8791) );
  CLKINVX1 U12292 ( .A(n8631), .Y(n8902) );
  OAI33X1 U12293 ( .A0(n1340), .A1(n187), .A2(n9741), .B0(n1461), .B1(n982), 
        .B2(n1339), .Y(n1459) );
  CLKMX2X2 U12294 ( .A(n8458), .B(n8459), .S0(n9136), .Y(n8552) );
  MX3XL U12295 ( .A(n8874), .B(n8866), .C(n8549), .S0(n8943), .S1(n8959), .Y(
        n8458) );
  MX3XL U12296 ( .A(n8826), .B(n8818), .C(n8548), .S0(n8941), .S1(n8958), .Y(
        n8459) );
  CLKMX2X2 U12297 ( .A(n8460), .B(n8461), .S0(n8923), .Y(n8572) );
  MX3XL U12298 ( .A(n8875), .B(n8867), .C(n8569), .S0(n8939), .S1(n8959), .Y(
        n8460) );
  MX3XL U12299 ( .A(n8827), .B(n8819), .C(n8568), .S0(n8941), .S1(n8959), .Y(
        n8461) );
  CLKMX2X2 U12300 ( .A(n8462), .B(n8463), .S0(n8923), .Y(n8592) );
  MX3XL U12301 ( .A(n8876), .B(n8868), .C(n8589), .S0(n8938), .S1(n8959), .Y(
        n8462) );
  MX3XL U12302 ( .A(n8828), .B(n8820), .C(n8588), .S0(n9140), .S1(n8959), .Y(
        n8463) );
  CLKMX2X2 U12303 ( .A(n8464), .B(n8465), .S0(n8920), .Y(n8612) );
  MX3XL U12304 ( .A(n8877), .B(n8869), .C(n8609), .S0(n8942), .S1(n8959), .Y(
        n8464) );
  MX3XL U12305 ( .A(n8829), .B(n8821), .C(n8608), .S0(n9140), .S1(n8959), .Y(
        n8465) );
  NAND2X1 U12306 ( .A(n9459), .B(n2453), .Y(n2415) );
  OAI33X1 U12307 ( .A0(n2290), .A1(n200), .A2(n9741), .B0(n2454), .B1(n9340), 
        .B2(n982), .Y(n2453) );
  NAND3X1 U12308 ( .A(N1656), .B(N1657), .C(n2585), .Y(n2454) );
  MX4X1 U12309 ( .A(\buff[4][2] ), .B(\buff[5][2] ), .C(\buff[6][2] ), .D(
        \buff[7][2] ), .S0(n9126), .S1(n9149), .Y(n9022) );
  MX4X1 U12310 ( .A(\buff[36][2] ), .B(\buff[37][2] ), .C(\buff[38][2] ), .D(
        \buff[39][2] ), .S0(n9133), .S1(n9149), .Y(n9012) );
  MX4X1 U12311 ( .A(\buff[4][3] ), .B(\buff[5][3] ), .C(\buff[6][3] ), .D(
        \buff[7][3] ), .S0(n9132), .S1(n9143), .Y(n9042) );
  MX4X1 U12312 ( .A(\buff[36][3] ), .B(\buff[37][3] ), .C(\buff[38][3] ), .D(
        \buff[39][3] ), .S0(n9132), .S1(n9142), .Y(n9032) );
  MX4X1 U12313 ( .A(\buff[36][4] ), .B(\buff[37][4] ), .C(\buff[38][4] ), .D(
        \buff[39][4] ), .S0(n9126), .S1(n9150), .Y(n9052) );
  MX4X1 U12314 ( .A(\buff[4][4] ), .B(\buff[5][4] ), .C(\buff[6][4] ), .D(
        \buff[7][4] ), .S0(n8919), .S1(n9151), .Y(n9062) );
  MX4X1 U12315 ( .A(\buff[4][5] ), .B(\buff[5][5] ), .C(\buff[6][5] ), .D(
        \buff[7][5] ), .S0(n9131), .S1(n9143), .Y(n9082) );
  MX4X1 U12316 ( .A(\buff[36][5] ), .B(\buff[37][5] ), .C(\buff[38][5] ), .D(
        \buff[39][5] ), .S0(n9127), .S1(n9151), .Y(n9072) );
  MX4X1 U12317 ( .A(\buff[20][2] ), .B(\buff[21][2] ), .C(\buff[22][2] ), .D(
        \buff[23][2] ), .S0(n9126), .S1(n9149), .Y(n9017) );
  MX4X1 U12318 ( .A(\buff[52][2] ), .B(\buff[53][2] ), .C(\buff[54][2] ), .D(
        \buff[55][2] ), .S0(n9133), .S1(n9148), .Y(n9007) );
  MX4X1 U12319 ( .A(n9018), .B(n9016), .C(n9017), .D(n9015), .S0(n9139), .S1(
        n8431), .Y(n9019) );
  MX4X1 U12320 ( .A(\buff[16][2] ), .B(\buff[17][2] ), .C(\buff[18][2] ), .D(
        \buff[19][2] ), .S0(n9127), .S1(n9149), .Y(n9018) );
  MX4X1 U12321 ( .A(\buff[24][2] ), .B(\buff[25][2] ), .C(\buff[26][2] ), .D(
        \buff[27][2] ), .S0(n9126), .S1(n9149), .Y(n9016) );
  MX4X1 U12322 ( .A(\buff[28][2] ), .B(\buff[29][2] ), .C(\buff[30][2] ), .D(
        \buff[31][2] ), .S0(n9127), .S1(n9149), .Y(n9015) );
  MX4X1 U12323 ( .A(\buff[20][3] ), .B(\buff[21][3] ), .C(\buff[22][3] ), .D(
        \buff[23][3] ), .S0(n9132), .S1(n8962), .Y(n9037) );
  MX4X1 U12324 ( .A(\buff[52][3] ), .B(\buff[53][3] ), .C(\buff[54][3] ), .D(
        \buff[55][3] ), .S0(n9127), .S1(n9147), .Y(n9027) );
  MX4X1 U12325 ( .A(n9038), .B(n9036), .C(n9037), .D(n9035), .S0(n9138), .S1(
        n9141), .Y(n9039) );
  MX4X1 U12326 ( .A(\buff[16][3] ), .B(\buff[17][3] ), .C(\buff[18][3] ), .D(
        \buff[19][3] ), .S0(n9132), .S1(n9144), .Y(n9038) );
  MX4X1 U12327 ( .A(\buff[24][3] ), .B(\buff[25][3] ), .C(\buff[26][3] ), .D(
        \buff[27][3] ), .S0(n9132), .S1(n8962), .Y(n9036) );
  MX4X1 U12328 ( .A(\buff[28][3] ), .B(\buff[29][3] ), .C(\buff[30][3] ), .D(
        \buff[31][3] ), .S0(n9132), .S1(n8961), .Y(n9035) );
  MX4X1 U12329 ( .A(\buff[20][4] ), .B(\buff[21][4] ), .C(\buff[22][4] ), .D(
        \buff[23][4] ), .S0(n9128), .S1(n9150), .Y(n9057) );
  MX4X1 U12330 ( .A(\buff[52][4] ), .B(\buff[53][4] ), .C(\buff[54][4] ), .D(
        \buff[55][4] ), .S0(n9128), .S1(n9150), .Y(n9047) );
  MX4X1 U12331 ( .A(n9058), .B(n9056), .C(n9057), .D(n9055), .S0(n8928), .S1(
        n9141), .Y(n9059) );
  MX4X1 U12332 ( .A(\buff[16][4] ), .B(\buff[17][4] ), .C(\buff[18][4] ), .D(
        \buff[19][4] ), .S0(n9128), .S1(n9150), .Y(n9058) );
  MX4X1 U12333 ( .A(\buff[24][4] ), .B(\buff[25][4] ), .C(\buff[26][4] ), .D(
        \buff[27][4] ), .S0(n9129), .S1(n9150), .Y(n9056) );
  MX4X1 U12334 ( .A(\buff[28][4] ), .B(\buff[29][4] ), .C(\buff[30][4] ), .D(
        \buff[31][4] ), .S0(n9128), .S1(n9150), .Y(n9055) );
  MX4X1 U12335 ( .A(\buff[20][5] ), .B(\buff[21][5] ), .C(\buff[22][5] ), .D(
        \buff[23][5] ), .S0(n8919), .S1(n9143), .Y(n9077) );
  MX4X1 U12336 ( .A(\buff[52][5] ), .B(\buff[53][5] ), .C(\buff[54][5] ), .D(
        \buff[55][5] ), .S0(n9125), .S1(n9151), .Y(n9067) );
  MX4X1 U12337 ( .A(n9078), .B(n9076), .C(n9077), .D(n9075), .S0(n8370), .S1(
        n9140), .Y(n9079) );
  MX4X1 U12338 ( .A(\buff[16][5] ), .B(\buff[17][5] ), .C(\buff[18][5] ), .D(
        \buff[19][5] ), .S0(n9131), .S1(n9146), .Y(n9078) );
  MX4X1 U12339 ( .A(\buff[24][5] ), .B(\buff[25][5] ), .C(\buff[26][5] ), .D(
        \buff[27][5] ), .S0(n9128), .S1(n9142), .Y(n9076) );
  MX4X1 U12340 ( .A(\buff[28][5] ), .B(\buff[29][5] ), .C(\buff[30][5] ), .D(
        \buff[31][5] ), .S0(n9129), .S1(n9151), .Y(n9075) );
  MX4X1 U12341 ( .A(\buff[0][1] ), .B(\buff[1][1] ), .C(\buff[2][1] ), .D(
        \buff[3][1] ), .S0(n9133), .S1(n9148), .Y(n9003) );
  MX4X1 U12342 ( .A(\buff[32][1] ), .B(\buff[33][1] ), .C(\buff[34][1] ), .D(
        \buff[35][1] ), .S0(n9134), .S1(n9147), .Y(n8993) );
  MX4X1 U12343 ( .A(\buff[48][2] ), .B(\buff[49][2] ), .C(\buff[50][2] ), .D(
        \buff[51][2] ), .S0(n9133), .S1(n9148), .Y(n9008) );
  MX4X1 U12344 ( .A(\buff[0][2] ), .B(\buff[1][2] ), .C(\buff[2][2] ), .D(
        \buff[3][2] ), .S0(n9126), .S1(n9149), .Y(n9023) );
  MX4X1 U12345 ( .A(\buff[32][2] ), .B(\buff[33][2] ), .C(\buff[34][2] ), .D(
        \buff[35][2] ), .S0(n9126), .S1(n9149), .Y(n9013) );
  MX4X1 U12346 ( .A(\buff[48][3] ), .B(\buff[49][3] ), .C(\buff[50][3] ), .D(
        \buff[51][3] ), .S0(n9126), .S1(n8955), .Y(n9028) );
  MX4X1 U12347 ( .A(\buff[0][3] ), .B(\buff[1][3] ), .C(\buff[2][3] ), .D(
        \buff[3][3] ), .S0(n9132), .S1(n9150), .Y(n9043) );
  MX4X1 U12348 ( .A(\buff[32][3] ), .B(\buff[33][3] ), .C(\buff[34][3] ), .D(
        \buff[35][3] ), .S0(n9132), .S1(n9144), .Y(n9033) );
  MX4X1 U12349 ( .A(\buff[48][4] ), .B(\buff[49][4] ), .C(\buff[50][4] ), .D(
        \buff[51][4] ), .S0(n9128), .S1(n9150), .Y(n9048) );
  MX4X1 U12350 ( .A(\buff[32][4] ), .B(\buff[33][4] ), .C(\buff[34][4] ), .D(
        \buff[35][4] ), .S0(n9128), .S1(n9150), .Y(n9053) );
  MX4X1 U12351 ( .A(\buff[0][4] ), .B(\buff[1][4] ), .C(\buff[2][4] ), .D(
        \buff[3][4] ), .S0(n8919), .S1(n9151), .Y(n9063) );
  MX4X1 U12352 ( .A(\buff[48][5] ), .B(\buff[49][5] ), .C(\buff[50][5] ), .D(
        \buff[51][5] ), .S0(n9129), .S1(n9151), .Y(n9068) );
  MX4X1 U12353 ( .A(\buff[0][5] ), .B(\buff[1][5] ), .C(\buff[2][5] ), .D(
        \buff[3][5] ), .S0(n9131), .S1(n9146), .Y(n9083) );
  MX4X1 U12354 ( .A(\buff[32][5] ), .B(\buff[33][5] ), .C(\buff[34][5] ), .D(
        \buff[35][5] ), .S0(n9126), .S1(n9151), .Y(n9073) );
  MX4X1 U12355 ( .A(\buff[12][2] ), .B(\buff[13][2] ), .C(\buff[14][2] ), .D(
        \buff[15][2] ), .S0(n9127), .S1(n9149), .Y(n9020) );
  MX4X1 U12356 ( .A(\buff[44][2] ), .B(\buff[45][2] ), .C(\buff[46][2] ), .D(
        \buff[47][2] ), .S0(n9133), .S1(n9148), .Y(n9010) );
  MX4X1 U12357 ( .A(\buff[12][3] ), .B(\buff[13][3] ), .C(\buff[14][3] ), .D(
        \buff[15][3] ), .S0(n9132), .S1(n8957), .Y(n9040) );
  MX4X1 U12358 ( .A(\buff[44][3] ), .B(\buff[45][3] ), .C(\buff[46][3] ), .D(
        \buff[47][3] ), .S0(n9132), .S1(n8957), .Y(n9030) );
  MX4X1 U12359 ( .A(\buff[44][4] ), .B(\buff[45][4] ), .C(\buff[46][4] ), .D(
        \buff[47][4] ), .S0(n9128), .S1(n9150), .Y(n9050) );
  MX4X1 U12360 ( .A(\buff[12][4] ), .B(\buff[13][4] ), .C(\buff[14][4] ), .D(
        \buff[15][4] ), .S0(n9126), .S1(n9151), .Y(n9060) );
  MX4X1 U12361 ( .A(\buff[12][5] ), .B(\buff[13][5] ), .C(\buff[14][5] ), .D(
        \buff[15][5] ), .S0(n9131), .S1(n9148), .Y(n9080) );
  MX4X1 U12362 ( .A(\buff[44][5] ), .B(\buff[45][5] ), .C(\buff[46][5] ), .D(
        \buff[47][5] ), .S0(n9128), .S1(n9151), .Y(n9070) );
  MX4X1 U12363 ( .A(\buff[60][2] ), .B(\buff[61][2] ), .C(\buff[62][2] ), .D(
        \buff[63][2] ), .S0(n9133), .S1(n9148), .Y(n9005) );
  MX4X1 U12364 ( .A(\buff[60][3] ), .B(\buff[61][3] ), .C(\buff[62][3] ), .D(
        \buff[63][3] ), .S0(n9127), .S1(n9149), .Y(n9025) );
  MX4X1 U12365 ( .A(\buff[60][4] ), .B(\buff[61][4] ), .C(\buff[62][4] ), .D(
        \buff[63][4] ), .S0(n9132), .S1(n9150), .Y(n9045) );
  MX4X1 U12366 ( .A(\buff[60][5] ), .B(\buff[61][5] ), .C(\buff[62][5] ), .D(
        \buff[63][5] ), .S0(n9127), .S1(n9151), .Y(n9065) );
  MX4X1 U12367 ( .A(\buff[8][1] ), .B(\buff[9][1] ), .C(\buff[10][1] ), .D(
        \buff[11][1] ), .S0(n9133), .S1(n9148), .Y(n9001) );
  MX4X1 U12368 ( .A(\buff[40][1] ), .B(\buff[41][1] ), .C(\buff[42][1] ), .D(
        \buff[43][1] ), .S0(n9134), .S1(n9147), .Y(n8991) );
  MX4X1 U12369 ( .A(\buff[8][2] ), .B(\buff[9][2] ), .C(\buff[10][2] ), .D(
        \buff[11][2] ), .S0(n9127), .S1(n9149), .Y(n9021) );
  MX4X1 U12370 ( .A(\buff[40][2] ), .B(\buff[41][2] ), .C(\buff[42][2] ), .D(
        \buff[43][2] ), .S0(n9133), .S1(n9149), .Y(n9011) );
  MX4X1 U12371 ( .A(\buff[8][3] ), .B(\buff[9][3] ), .C(\buff[10][3] ), .D(
        \buff[11][3] ), .S0(n9132), .S1(n9152), .Y(n9041) );
  MX4X1 U12372 ( .A(\buff[40][3] ), .B(\buff[41][3] ), .C(\buff[42][3] ), .D(
        \buff[43][3] ), .S0(n9132), .S1(n8955), .Y(n9031) );
  MX4X1 U12373 ( .A(\buff[40][4] ), .B(\buff[41][4] ), .C(\buff[42][4] ), .D(
        \buff[43][4] ), .S0(n9129), .S1(n9150), .Y(n9051) );
  MX4X1 U12374 ( .A(\buff[8][4] ), .B(\buff[9][4] ), .C(\buff[10][4] ), .D(
        \buff[11][4] ), .S0(n9129), .S1(n9151), .Y(n9061) );
  MX4X1 U12375 ( .A(\buff[8][5] ), .B(\buff[9][5] ), .C(\buff[10][5] ), .D(
        \buff[11][5] ), .S0(n9131), .S1(n9143), .Y(n9081) );
  MX4X1 U12376 ( .A(\buff[40][5] ), .B(\buff[41][5] ), .C(\buff[42][5] ), .D(
        \buff[43][5] ), .S0(n9129), .S1(n9151), .Y(n9071) );
  MX4X1 U12377 ( .A(\buff[56][2] ), .B(\buff[57][2] ), .C(\buff[58][2] ), .D(
        \buff[59][2] ), .S0(n9133), .S1(n9148), .Y(n9006) );
  MX4X1 U12378 ( .A(\buff[56][3] ), .B(\buff[57][3] ), .C(\buff[58][3] ), .D(
        \buff[59][3] ), .S0(n9126), .S1(n9149), .Y(n9026) );
  MX4X1 U12379 ( .A(\buff[56][4] ), .B(\buff[57][4] ), .C(\buff[58][4] ), .D(
        \buff[59][4] ), .S0(n9129), .S1(n9150), .Y(n9046) );
  MX4X1 U12380 ( .A(\buff[56][5] ), .B(\buff[57][5] ), .C(\buff[58][5] ), .D(
        \buff[59][5] ), .S0(n9129), .S1(n9151), .Y(n9066) );
  CLKINVX1 U12381 ( .A(cmd_valid), .Y(n9717) );
  MXI3X1 U12382 ( .A(n8858), .B(n8850), .C(n8543), .S0(n8942), .S1(n8959), .Y(
        n8542) );
  CLKINVX1 U12383 ( .A(\buff[19][3] ), .Y(n8850) );
  CLKINVX1 U12384 ( .A(\buff[15][3] ), .Y(n8858) );
  MXI3X1 U12385 ( .A(n8859), .B(n8851), .C(n8563), .S0(n8938), .S1(n8959), .Y(
        n8562) );
  CLKINVX1 U12386 ( .A(\buff[19][4] ), .Y(n8851) );
  CLKINVX1 U12387 ( .A(\buff[15][4] ), .Y(n8859) );
  MXI3X1 U12388 ( .A(n8860), .B(n8852), .C(n8583), .S0(n8942), .S1(n8959), .Y(
        n8582) );
  CLKINVX1 U12389 ( .A(\buff[19][5] ), .Y(n8852) );
  CLKINVX1 U12390 ( .A(\buff[15][5] ), .Y(n8860) );
  MXI3X1 U12391 ( .A(n8861), .B(n8853), .C(n8603), .S0(n8939), .S1(n8959), .Y(
        n8602) );
  CLKINVX1 U12392 ( .A(\buff[19][6] ), .Y(n8853) );
  CLKINVX1 U12393 ( .A(\buff[15][6] ), .Y(n8861) );
  MXI3X1 U12394 ( .A(n8862), .B(n8854), .C(n8623), .S0(n8942), .S1(n8959), .Y(
        n8622) );
  CLKINVX1 U12395 ( .A(\buff[15][7] ), .Y(n8862) );
  CLKINVX1 U12396 ( .A(\buff[19][7] ), .Y(n8854) );
  CLKINVX1 U12397 ( .A(\buff[3][0] ), .Y(n8879) );
  CLKINVX1 U12398 ( .A(\buff[3][1] ), .Y(n8880) );
  MX4X1 U12399 ( .A(\buff[24][2] ), .B(\buff[28][2] ), .C(\buff[26][2] ), .D(
        \buff[30][2] ), .S0(n8944), .S1(n8960), .Y(n8466) );
  MX4X1 U12400 ( .A(\buff[24][3] ), .B(\buff[28][3] ), .C(\buff[26][3] ), .D(
        \buff[30][3] ), .S0(n8945), .S1(n8960), .Y(n8467) );
  MX4X1 U12401 ( .A(\buff[24][4] ), .B(\buff[28][4] ), .C(\buff[26][4] ), .D(
        \buff[30][4] ), .S0(n8942), .S1(n8960), .Y(n8468) );
  MX4X1 U12402 ( .A(\buff[24][5] ), .B(\buff[28][5] ), .C(\buff[26][5] ), .D(
        \buff[30][5] ), .S0(n8935), .S1(n8959), .Y(n8469) );
  MX4X1 U12403 ( .A(\buff[24][6] ), .B(\buff[28][6] ), .C(\buff[26][6] ), .D(
        \buff[30][6] ), .S0(n8953), .S1(n8959), .Y(n8470) );
  CLKINVX1 U12404 ( .A(\buff[43][0] ), .Y(n8815) );
  CLKINVX1 U12405 ( .A(\buff[51][0] ), .Y(n8799) );
  CLKINVX1 U12406 ( .A(\buff[35][0] ), .Y(n8831) );
  CLKINVX1 U12407 ( .A(\buff[43][1] ), .Y(n8816) );
  CLKINVX1 U12408 ( .A(\buff[11][1] ), .Y(n8864) );
  CLKINVX1 U12409 ( .A(\buff[51][1] ), .Y(n8800) );
  CLKINVX1 U12410 ( .A(\buff[35][1] ), .Y(n8832) );
  CLKINVX1 U12411 ( .A(\buff[39][0] ), .Y(n8823) );
  CLKINVX1 U12412 ( .A(\buff[7][0] ), .Y(n8871) );
  CLKINVX1 U12413 ( .A(\buff[47][0] ), .Y(n8807) );
  CLKINVX1 U12414 ( .A(\buff[31][0] ), .Y(n8839) );
  CLKINVX1 U12415 ( .A(\buff[39][1] ), .Y(n8824) );
  CLKINVX1 U12416 ( .A(\buff[47][1] ), .Y(n8808) );
  CLKINVX1 U12417 ( .A(\buff[31][1] ), .Y(n8840) );
  MXI4X1 U12418 ( .A(n8529), .B(n8667), .C(n8528), .D(n8668), .S0(n8962), .S1(
        n8921), .Y(n8666) );
  MXI2X1 U12419 ( .A(\buff[43][2] ), .B(\buff[47][2] ), .S0(n8930), .Y(n8668)
         );
  MXI2X1 U12420 ( .A(\buff[11][2] ), .B(\buff[15][2] ), .S0(n8939), .Y(n8667)
         );
  MXI4X1 U12421 ( .A(n8549), .B(n8680), .C(n8548), .D(n8681), .S0(n8961), .S1(
        n8921), .Y(n8679) );
  MXI2X1 U12422 ( .A(\buff[43][3] ), .B(\buff[47][3] ), .S0(n8943), .Y(n8681)
         );
  MXI2X1 U12423 ( .A(\buff[11][3] ), .B(\buff[15][3] ), .S0(n8943), .Y(n8680)
         );
  MXI4X1 U12424 ( .A(n8569), .B(n8693), .C(n8568), .D(n8694), .S0(n8962), .S1(
        n8922), .Y(n8692) );
  MXI2X1 U12425 ( .A(\buff[43][4] ), .B(\buff[47][4] ), .S0(n8944), .Y(n8694)
         );
  MXI2X1 U12426 ( .A(\buff[11][4] ), .B(\buff[15][4] ), .S0(n8944), .Y(n8693)
         );
  MXI4X1 U12427 ( .A(n8589), .B(n8706), .C(n8588), .D(n8707), .S0(n8962), .S1(
        n8922), .Y(n8705) );
  MXI2X1 U12428 ( .A(\buff[43][5] ), .B(\buff[47][5] ), .S0(n8937), .Y(n8707)
         );
  MXI2X1 U12429 ( .A(\buff[11][5] ), .B(\buff[15][5] ), .S0(n8940), .Y(n8706)
         );
  MXI4X1 U12430 ( .A(n8609), .B(n8719), .C(n8608), .D(n8720), .S0(n8961), .S1(
        n8922), .Y(n8718) );
  MXI2X1 U12431 ( .A(\buff[43][6] ), .B(\buff[47][6] ), .S0(n8945), .Y(n8720)
         );
  MXI2X1 U12432 ( .A(\buff[11][6] ), .B(\buff[15][6] ), .S0(n8940), .Y(n8719)
         );
  MXI4X1 U12433 ( .A(n8523), .B(n8661), .C(n8521), .D(n8662), .S0(n8961), .S1(
        n8921), .Y(n8660) );
  MXI2X1 U12434 ( .A(\buff[51][2] ), .B(\buff[55][2] ), .S0(n8943), .Y(n8662)
         );
  MXI2X1 U12435 ( .A(\buff[19][2] ), .B(\buff[23][2] ), .S0(n8943), .Y(n8661)
         );
  MXI4X1 U12436 ( .A(n8543), .B(n8674), .C(n8541), .D(n8675), .S0(n8961), .S1(
        n8921), .Y(n8673) );
  MXI2X1 U12437 ( .A(\buff[51][3] ), .B(\buff[55][3] ), .S0(n8938), .Y(n8675)
         );
  MXI2X1 U12438 ( .A(\buff[19][3] ), .B(\buff[23][3] ), .S0(n8938), .Y(n8674)
         );
  MXI4X1 U12439 ( .A(n8563), .B(n8687), .C(n8561), .D(n8688), .S0(n8962), .S1(
        n8921), .Y(n8686) );
  MXI2X1 U12440 ( .A(\buff[51][4] ), .B(\buff[55][4] ), .S0(n8943), .Y(n8688)
         );
  MXI2X1 U12441 ( .A(\buff[19][4] ), .B(\buff[23][4] ), .S0(n8943), .Y(n8687)
         );
  MXI4X1 U12442 ( .A(n8583), .B(n8700), .C(n8581), .D(n8701), .S0(n8961), .S1(
        n8922), .Y(n8699) );
  MXI2X1 U12443 ( .A(\buff[51][5] ), .B(\buff[55][5] ), .S0(n8944), .Y(n8701)
         );
  MXI2X1 U12444 ( .A(\buff[19][5] ), .B(\buff[23][5] ), .S0(n8944), .Y(n8700)
         );
  MXI4X1 U12445 ( .A(n8603), .B(n8713), .C(n8601), .D(n8714), .S0(n8961), .S1(
        n8922), .Y(n8712) );
  MXI2X1 U12446 ( .A(\buff[51][6] ), .B(\buff[55][6] ), .S0(n9140), .Y(n8714)
         );
  MXI2X1 U12447 ( .A(\buff[19][6] ), .B(\buff[23][6] ), .S0(n9140), .Y(n8713)
         );
  MXI4X1 U12448 ( .A(n8527), .B(n8664), .C(n8525), .D(n8665), .S0(n8961), .S1(
        n8921), .Y(n8663) );
  MXI2X1 U12449 ( .A(\buff[35][2] ), .B(\buff[39][2] ), .S0(n8943), .Y(n8665)
         );
  MXI2X1 U12450 ( .A(\buff[3][2] ), .B(\buff[7][2] ), .S0(n8943), .Y(n8664) );
  MXI4X1 U12451 ( .A(n8547), .B(n8677), .C(n8545), .D(n8678), .S0(n8962), .S1(
        n8921), .Y(n8676) );
  MXI2X1 U12452 ( .A(\buff[35][3] ), .B(\buff[39][3] ), .S0(n8949), .Y(n8678)
         );
  MXI2X1 U12453 ( .A(\buff[3][3] ), .B(\buff[7][3] ), .S0(n8953), .Y(n8677) );
  MXI4X1 U12454 ( .A(n8567), .B(n8690), .C(n8565), .D(n8691), .S0(n8961), .S1(
        n8921), .Y(n8689) );
  MXI2X1 U12455 ( .A(\buff[35][4] ), .B(\buff[39][4] ), .S0(n8943), .Y(n8691)
         );
  MXI2X1 U12456 ( .A(\buff[3][4] ), .B(\buff[7][4] ), .S0(n8943), .Y(n8690) );
  MXI4X1 U12457 ( .A(n8587), .B(n8703), .C(n8585), .D(n8704), .S0(n8961), .S1(
        n8922), .Y(n8702) );
  MXI2X1 U12458 ( .A(\buff[35][5] ), .B(\buff[39][5] ), .S0(n8944), .Y(n8704)
         );
  MXI2X1 U12459 ( .A(\buff[3][5] ), .B(\buff[7][5] ), .S0(n8945), .Y(n8703) );
  MXI4X1 U12460 ( .A(n8607), .B(n8716), .C(n8605), .D(n8717), .S0(n8962), .S1(
        n8922), .Y(n8715) );
  MXI2X1 U12461 ( .A(\buff[35][6] ), .B(\buff[39][6] ), .S0(n8937), .Y(n8717)
         );
  MXI2X1 U12462 ( .A(\buff[3][6] ), .B(\buff[7][6] ), .S0(n8938), .Y(n8716) );
  MX4X1 U12463 ( .A(\buff[48][4] ), .B(\buff[52][4] ), .C(\buff[50][4] ), .D(
        \buff[54][4] ), .S0(n8951), .S1(n9142), .Y(n8554) );
  MX4X1 U12464 ( .A(\buff[32][4] ), .B(\buff[36][4] ), .C(\buff[34][4] ), .D(
        \buff[38][4] ), .S0(n8950), .S1(n9143), .Y(n8556) );
  MX4X1 U12465 ( .A(\buff[48][5] ), .B(\buff[52][5] ), .C(\buff[50][5] ), .D(
        \buff[54][5] ), .S0(n8950), .S1(n9151), .Y(n8574) );
  MX4X1 U12466 ( .A(\buff[32][5] ), .B(\buff[36][5] ), .C(\buff[34][5] ), .D(
        \buff[38][5] ), .S0(n8950), .S1(n9146), .Y(n8576) );
  MX4X1 U12467 ( .A(\buff[48][6] ), .B(\buff[52][6] ), .C(\buff[50][6] ), .D(
        \buff[54][6] ), .S0(n8950), .S1(n8956), .Y(n8594) );
  MX4X1 U12468 ( .A(\buff[32][6] ), .B(\buff[36][6] ), .C(\buff[34][6] ), .D(
        \buff[38][6] ), .S0(n8950), .S1(n9143), .Y(n8596) );
  MX4X1 U12469 ( .A(\buff[48][7] ), .B(\buff[52][7] ), .C(\buff[50][7] ), .D(
        \buff[54][7] ), .S0(n8949), .S1(n8964), .Y(n8614) );
  MX4X1 U12470 ( .A(\buff[32][7] ), .B(\buff[36][7] ), .C(\buff[34][7] ), .D(
        \buff[38][7] ), .S0(n8949), .S1(n8956), .Y(n8616) );
  OAI21XL U12471 ( .A0(n2581), .A1(n9340), .B0(n9744), .Y(n2567) );
  NOR3XL U12472 ( .A(IROM_A[0]), .B(IROM_A[2]), .C(IROM_A[1]), .Y(n2568) );
  MXI2X1 U12473 ( .A(\buff[1][7] ), .B(\buff[5][7] ), .S0(n8945), .Y(n8627) );
  CLKMX2X2 U12474 ( .A(n8471), .B(n8472), .S0(n8920), .Y(n8632) );
  MX3XL U12475 ( .A(n8878), .B(n8870), .C(n8629), .S0(n8942), .S1(n8958), .Y(
        n8471) );
  MX3XL U12476 ( .A(n8830), .B(n8822), .C(n8628), .S0(n8942), .S1(n8959), .Y(
        n8472) );
  MXI2X1 U12477 ( .A(\buff[41][7] ), .B(\buff[45][7] ), .S0(n8945), .Y(n8628)
         );
  MXI2X1 U12478 ( .A(\buff[9][7] ), .B(\buff[13][7] ), .S0(n8945), .Y(n8629)
         );
  OAI2BB2XL U12479 ( .B0(n8385), .B1(n2565), .A0N(N1748), .A1N(n2566), .Y(
        n3113) );
  OAI2BB2XL U12480 ( .B0(n8383), .B1(n2565), .A0N(N1747), .A1N(n2566), .Y(
        n3114) );
  OAI2BB2XL U12481 ( .B0(n2584), .B1(n2565), .A0N(N1746), .A1N(n2566), .Y(
        n3115) );
  OAI2BB2XL U12482 ( .B0(n2585), .B1(n2565), .A0N(N1745), .A1N(n2566), .Y(
        n3116) );
  OAI2BB2XL U12483 ( .B0(n2581), .B1(n2565), .A0N(N1749), .A1N(n2566), .Y(
        n3119) );
  MXI2X1 U12484 ( .A(\buff[27][6] ), .B(\buff[31][6] ), .S0(n8939), .Y(n8723)
         );
  MXI2X1 U12485 ( .A(\buff[27][7] ), .B(\buff[31][7] ), .S0(n8946), .Y(n8736)
         );
  MXI2X1 U12486 ( .A(n8473), .B(n8787), .S0(n9136), .Y(n8790) );
  MX4X1 U12487 ( .A(\buff[56][7] ), .B(\buff[60][7] ), .C(\buff[58][7] ), .D(
        \buff[62][7] ), .S0(n8948), .S1(n8960), .Y(n8787) );
  MX4X1 U12488 ( .A(\buff[4][6] ), .B(\buff[5][6] ), .C(\buff[6][6] ), .D(
        \buff[7][6] ), .S0(n9130), .S1(n9144), .Y(n9102) );
  MX4X1 U12489 ( .A(\buff[36][6] ), .B(\buff[37][6] ), .C(\buff[38][6] ), .D(
        \buff[39][6] ), .S0(n9131), .S1(n9151), .Y(n9092) );
  MX4X1 U12490 ( .A(n9098), .B(n9096), .C(n9097), .D(n9095), .S0(n9511), .S1(
        n8431), .Y(n9099) );
  MX4X1 U12491 ( .A(\buff[16][6] ), .B(\buff[17][6] ), .C(\buff[18][6] ), .D(
        \buff[19][6] ), .S0(n9130), .S1(n9142), .Y(n9098) );
  MX4X1 U12492 ( .A(\buff[24][6] ), .B(\buff[25][6] ), .C(\buff[26][6] ), .D(
        \buff[27][6] ), .S0(n9130), .S1(n9142), .Y(n9096) );
  MX4X1 U12493 ( .A(\buff[28][6] ), .B(\buff[29][6] ), .C(\buff[30][6] ), .D(
        \buff[31][6] ), .S0(n9130), .S1(n9149), .Y(n9095) );
  MX4X1 U12494 ( .A(\buff[4][7] ), .B(\buff[5][7] ), .C(\buff[6][7] ), .D(
        \buff[7][7] ), .S0(n9517), .S1(n9149), .Y(n9122) );
  MX4X1 U12495 ( .A(\buff[36][7] ), .B(\buff[37][7] ), .C(\buff[38][7] ), .D(
        \buff[39][7] ), .S0(n9129), .S1(n9143), .Y(n9112) );
  MX4X1 U12496 ( .A(n9118), .B(n9116), .C(n9117), .D(n9115), .S0(n9511), .S1(
        n9140), .Y(n9119) );
  MX4X1 U12497 ( .A(\buff[16][7] ), .B(\buff[17][7] ), .C(\buff[18][7] ), .D(
        \buff[19][7] ), .S0(n9517), .S1(n9142), .Y(n9118) );
  MX4X1 U12498 ( .A(\buff[24][7] ), .B(\buff[25][7] ), .C(\buff[26][7] ), .D(
        \buff[27][7] ), .S0(n9129), .S1(n9142), .Y(n9116) );
  MX4X1 U12499 ( .A(\buff[28][7] ), .B(\buff[29][7] ), .C(\buff[30][7] ), .D(
        \buff[31][7] ), .S0(n9517), .S1(n9142), .Y(n9115) );
  MX4X1 U12500 ( .A(\buff[20][6] ), .B(\buff[21][6] ), .C(\buff[22][6] ), .D(
        \buff[23][6] ), .S0(n9130), .S1(n8959), .Y(n9097) );
  MX4X1 U12501 ( .A(\buff[52][6] ), .B(\buff[53][6] ), .C(\buff[54][6] ), .D(
        \buff[55][6] ), .S0(n9131), .S1(n8961), .Y(n9087) );
  MX4X1 U12502 ( .A(\buff[52][7] ), .B(\buff[53][7] ), .C(\buff[54][7] ), .D(
        \buff[55][7] ), .S0(n9130), .S1(n9146), .Y(n9107) );
  MX4X1 U12503 ( .A(\buff[20][7] ), .B(\buff[21][7] ), .C(\buff[22][7] ), .D(
        \buff[23][7] ), .S0(n9517), .S1(n9150), .Y(n9117) );
  MX4X1 U12504 ( .A(\buff[48][6] ), .B(\buff[49][6] ), .C(\buff[50][6] ), .D(
        \buff[51][6] ), .S0(n9131), .S1(n8955), .Y(n9088) );
  MX4X1 U12505 ( .A(\buff[0][6] ), .B(\buff[1][6] ), .C(\buff[2][6] ), .D(
        \buff[3][6] ), .S0(n9130), .S1(n9148), .Y(n9103) );
  MX4X1 U12506 ( .A(\buff[32][6] ), .B(\buff[33][6] ), .C(\buff[34][6] ), .D(
        \buff[35][6] ), .S0(n9131), .S1(n9149), .Y(n9093) );
  MX4X1 U12507 ( .A(\buff[48][7] ), .B(\buff[49][7] ), .C(\buff[50][7] ), .D(
        \buff[51][7] ), .S0(n9130), .S1(n9142), .Y(n9108) );
  MX4X1 U12508 ( .A(\buff[0][7] ), .B(\buff[1][7] ), .C(\buff[2][7] ), .D(
        \buff[3][7] ), .S0(n9517), .S1(n9143), .Y(n9123) );
  MX4X1 U12509 ( .A(\buff[32][7] ), .B(\buff[33][7] ), .C(\buff[34][7] ), .D(
        \buff[35][7] ), .S0(n9128), .S1(n9142), .Y(n9113) );
  MX4X1 U12510 ( .A(\buff[12][6] ), .B(\buff[13][6] ), .C(\buff[14][6] ), .D(
        \buff[15][6] ), .S0(n9130), .S1(n9151), .Y(n9100) );
  MX4X1 U12511 ( .A(\buff[44][6] ), .B(\buff[45][6] ), .C(\buff[46][6] ), .D(
        \buff[47][6] ), .S0(n9131), .S1(n8962), .Y(n9090) );
  MX4X1 U12512 ( .A(\buff[12][7] ), .B(\buff[13][7] ), .C(\buff[14][7] ), .D(
        \buff[15][7] ), .S0(n8373), .S1(n9142), .Y(n9120) );
  MX4X1 U12513 ( .A(\buff[44][7] ), .B(\buff[45][7] ), .C(\buff[46][7] ), .D(
        \buff[47][7] ), .S0(n9130), .S1(n9143), .Y(n9110) );
  MX4X1 U12514 ( .A(\buff[60][6] ), .B(\buff[61][6] ), .C(\buff[62][6] ), .D(
        \buff[63][6] ), .S0(n9131), .S1(n9146), .Y(n9085) );
  MX4X1 U12515 ( .A(\buff[60][7] ), .B(\buff[61][7] ), .C(\buff[62][7] ), .D(
        \buff[63][7] ), .S0(n9130), .S1(n9149), .Y(n9105) );
  MX4X1 U12516 ( .A(\buff[8][6] ), .B(\buff[9][6] ), .C(\buff[10][6] ), .D(
        \buff[11][6] ), .S0(n9130), .S1(n9150), .Y(n9101) );
  MX4X1 U12517 ( .A(\buff[40][6] ), .B(\buff[41][6] ), .C(\buff[42][6] ), .D(
        \buff[43][6] ), .S0(n9131), .S1(n9145), .Y(n9091) );
  MX4X1 U12518 ( .A(\buff[8][7] ), .B(\buff[9][7] ), .C(\buff[10][7] ), .D(
        \buff[11][7] ), .S0(n9128), .S1(n9143), .Y(n9121) );
  MX4X1 U12519 ( .A(\buff[40][7] ), .B(\buff[41][7] ), .C(\buff[42][7] ), .D(
        \buff[43][7] ), .S0(n8919), .S1(n9142), .Y(n9111) );
  MX4X1 U12520 ( .A(\buff[56][6] ), .B(\buff[57][6] ), .C(\buff[58][6] ), .D(
        \buff[59][6] ), .S0(n9131), .S1(n9143), .Y(n9086) );
  MX4X1 U12521 ( .A(\buff[56][7] ), .B(\buff[57][7] ), .C(\buff[58][7] ), .D(
        \buff[59][7] ), .S0(n9130), .S1(n9150), .Y(n9106) );
  CLKINVX1 U12522 ( .A(\buff[3][2] ), .Y(n8881) );
  CLKINVX1 U12523 ( .A(\buff[3][3] ), .Y(n8882) );
  CLKINVX1 U12524 ( .A(\buff[3][4] ), .Y(n8883) );
  CLKINVX1 U12525 ( .A(\buff[3][5] ), .Y(n8884) );
  MX4X1 U12526 ( .A(\buff[24][7] ), .B(\buff[28][7] ), .C(\buff[26][7] ), .D(
        \buff[30][7] ), .S0(n8938), .S1(n8959), .Y(n8473) );
  CLKINVX1 U12527 ( .A(\buff[43][2] ), .Y(n8817) );
  CLKINVX1 U12528 ( .A(\buff[51][2] ), .Y(n8801) );
  CLKINVX1 U12529 ( .A(\buff[35][2] ), .Y(n8833) );
  CLKINVX1 U12530 ( .A(\buff[43][3] ), .Y(n8818) );
  CLKINVX1 U12531 ( .A(\buff[51][3] ), .Y(n8802) );
  CLKINVX1 U12532 ( .A(\buff[35][3] ), .Y(n8834) );
  CLKINVX1 U12533 ( .A(\buff[43][4] ), .Y(n8819) );
  CLKINVX1 U12534 ( .A(\buff[51][4] ), .Y(n8803) );
  CLKINVX1 U12535 ( .A(\buff[35][4] ), .Y(n8835) );
  CLKINVX1 U12536 ( .A(\buff[43][5] ), .Y(n8820) );
  CLKINVX1 U12537 ( .A(\buff[51][5] ), .Y(n8804) );
  CLKINVX1 U12538 ( .A(\buff[35][5] ), .Y(n8836) );
  CLKINVX1 U12539 ( .A(\buff[43][6] ), .Y(n8821) );
  CLKINVX1 U12540 ( .A(\buff[51][6] ), .Y(n8805) );
  CLKINVX1 U12541 ( .A(\buff[35][6] ), .Y(n8837) );
  CLKINVX1 U12542 ( .A(\buff[39][2] ), .Y(n8825) );
  CLKINVX1 U12543 ( .A(\buff[7][2] ), .Y(n8873) );
  CLKINVX1 U12544 ( .A(\buff[47][2] ), .Y(n8809) );
  CLKINVX1 U12545 ( .A(\buff[31][2] ), .Y(n8841) );
  CLKINVX1 U12546 ( .A(\buff[39][3] ), .Y(n8826) );
  CLKINVX1 U12547 ( .A(\buff[7][3] ), .Y(n8874) );
  CLKINVX1 U12548 ( .A(\buff[47][3] ), .Y(n8810) );
  CLKINVX1 U12549 ( .A(\buff[31][3] ), .Y(n8842) );
  CLKINVX1 U12550 ( .A(\buff[39][4] ), .Y(n8827) );
  CLKINVX1 U12551 ( .A(\buff[7][4] ), .Y(n8875) );
  CLKINVX1 U12552 ( .A(\buff[47][4] ), .Y(n8811) );
  CLKINVX1 U12553 ( .A(\buff[31][4] ), .Y(n8843) );
  CLKINVX1 U12554 ( .A(\buff[39][5] ), .Y(n8828) );
  CLKINVX1 U12555 ( .A(\buff[7][5] ), .Y(n8876) );
  CLKINVX1 U12556 ( .A(\buff[47][5] ), .Y(n8812) );
  CLKINVX1 U12557 ( .A(\buff[31][5] ), .Y(n8844) );
  CLKINVX1 U12558 ( .A(\buff[39][6] ), .Y(n8829) );
  CLKINVX1 U12559 ( .A(\buff[7][6] ), .Y(n8877) );
  CLKINVX1 U12560 ( .A(\buff[47][6] ), .Y(n8813) );
  CLKINVX1 U12561 ( .A(\buff[31][6] ), .Y(n8845) );
  MXI4X1 U12562 ( .A(n8629), .B(n8732), .C(n8628), .D(n8733), .S0(n8962), .S1(
        n8922), .Y(n8731) );
  MXI2X1 U12563 ( .A(\buff[43][7] ), .B(\buff[47][7] ), .S0(n9140), .Y(n8733)
         );
  MXI2X1 U12564 ( .A(\buff[11][7] ), .B(\buff[15][7] ), .S0(n8948), .Y(n8732)
         );
  MXI4X1 U12565 ( .A(n8623), .B(n8726), .C(n8621), .D(n8727), .S0(n8962), .S1(
        n8922), .Y(n8725) );
  MXI2X1 U12566 ( .A(\buff[51][7] ), .B(\buff[55][7] ), .S0(n8946), .Y(n8727)
         );
  MXI2X1 U12567 ( .A(\buff[19][7] ), .B(\buff[23][7] ), .S0(n8946), .Y(n8726)
         );
  MXI4X1 U12568 ( .A(n8627), .B(n8729), .C(n8625), .D(n8730), .S0(n8962), .S1(
        n8922), .Y(n8728) );
  MXI2X1 U12569 ( .A(\buff[35][7] ), .B(\buff[39][7] ), .S0(n8946), .Y(n8730)
         );
  MXI2X1 U12570 ( .A(\buff[3][7] ), .B(\buff[7][7] ), .S0(n8946), .Y(n8729) );
  NOR3X1 U12571 ( .A(n2590), .B(n2589), .C(n2591), .Y(n292) );
  CLKINVX1 U12572 ( .A(\buff[3][6] ), .Y(n8885) );
  CLKINVX1 U12573 ( .A(\buff[3][7] ), .Y(n8886) );
  CLKBUFX3 U12574 ( .A(n2502), .Y(n9348) );
  NOR3X1 U12575 ( .A(n2591), .B(n2589), .C(n9748), .Y(n2502) );
  CLKINVX1 U12576 ( .A(\buff[43][7] ), .Y(n8822) );
  CLKINVX1 U12577 ( .A(\buff[11][7] ), .Y(n8870) );
  CLKINVX1 U12578 ( .A(\buff[51][7] ), .Y(n8806) );
  CLKINVX1 U12579 ( .A(\buff[35][7] ), .Y(n8838) );
  CLKINVX1 U12580 ( .A(\buff[39][7] ), .Y(n8830) );
  CLKINVX1 U12581 ( .A(\buff[47][7] ), .Y(n8814) );
  CLKINVX1 U12582 ( .A(\buff[31][7] ), .Y(n8846) );
  CLKBUFX3 U12583 ( .A(n293), .Y(n9606) );
  NOR3X1 U12584 ( .A(n2590), .B(n2589), .C(n9738), .Y(n293) );
  NAND3X2 U12585 ( .A(n2584), .B(N1661), .C(n8383), .Y(n1024) );
  NAND3X2 U12586 ( .A(N1659), .B(N1661), .C(n8383), .Y(n704) );
  NAND3X2 U12587 ( .A(n8383), .B(N1659), .C(n8385), .Y(n1974) );
  NAND3X2 U12588 ( .A(n8393), .B(N1661), .C(n7474), .Y(n365) );
  NAND3X2 U12589 ( .A(N1659), .B(n8393), .C(n8385), .Y(n1339) );
  AOI2BB2X1 U12590 ( .B0(n8373), .B1(n2552), .A0N(n9740), .A1N(n8373), .Y(
        n2550) );
  NAND3X1 U12591 ( .A(n2586), .B(n2587), .C(n2585), .Y(n981) );
  NOR3X1 U12592 ( .A(n9748), .B(n2591), .C(n9747), .Y(n2546) );
  NOR3X1 U12593 ( .A(n2591), .B(n2590), .C(n9747), .Y(n2557) );
  NAND3X1 U12594 ( .A(n8383), .B(n2584), .C(n8385), .Y(n2289) );
  OR4X1 U12595 ( .A(n8393), .B(N1659), .C(\cnt[6] ), .D(N1661), .Y(n9667) );
  OR4X1 U12596 ( .A(N1658), .B(N1657), .C(n9317), .D(n9667), .Y(N1677) );
endmodule

